* File: Coin_bank.pex.sp
* Created: Sun Jan 14 15:06:01 2024
* Program "Calibre xRC"
* Version "v2021.3_35.19"
* 
.include "Coin_bank.pex.sp.pex"
.subckt COIN_BANK  State1 State0 S3 S2 S1 S0 Mo3 Mo2 Mo1 Mo0 Init3 Init2 Init1 Init0 M3 M2 M1 M0 Store Power Clk VDD VSS
* 
* M3	M3
* M2	M2
* M1	M1
* M0	M0
* CLK	CLK
* VSS	VSS
* VDD	VDD
* MO3	MO3
* MO2	MO2
* MO1	MO1
* S0	S0
* POWER	POWER
* MO0	MO0
* S2	S2
* STATE1	STATE1
* STATE0	STATE0
* STORE	STORE
* S1	S1
* S3	S3
* INIT3	INIT3
* INIT2	INIT2
* INIT1	INIT1
* INIT0	INIT0
mX0/X0/M0 N_X0/X0/6_X0/X0/M0_d N_9_X0/X0/M0_g N_VSS_X0/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX0/X0/M1 N_47_X0/X0/M1_d N_10_X0/X0/M1_g N_X0/X0/6_X0/X0/M1_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX0/X0/M2 N_47_X0/X0/M2_d N_9_X0/X0/M2_g N_VDD_X0/X0/M2_s N_VDD_X0/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX0/X0/M3 N_VDD_X0/X0/M3_d N_10_X0/X0/M3_g N_47_X0/X0/M3_s N_VDD_X0/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX0/X1/M0 N_11_X0/X1/M0_d N_47_X0/X1/M0_g N_VSS_X0/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX0/X1/M1 N_11_X0/X1/M1_d N_47_X0/X1/M1_g N_VDD_X0/X1/M1_s N_VDD_X0/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX1/X0/M0 N_X1/X0/6_X1/X0/M0_d N_STATE1_X1/X0/M0_g N_VSS_X1/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX1/X0/M1 N_48_X1/X0/M1_d N_STATE0_X1/X0/M1_g N_X1/X0/6_X1/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX1/X0/M2 N_48_X1/X0/M2_d N_STATE1_X1/X0/M2_g N_VDD_X1/X0/M2_s N_VDD_X1/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX1/X0/M3 N_VDD_X1/X0/M3_d N_STATE0_X1/X0/M3_g N_48_X1/X0/M3_s N_VDD_X1/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX1/X1/M0 N_S3_X1/X1/M0_d N_48_X1/X1/M0_g N_VSS_X1/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX1/X1/M1 N_S3_X1/X1/M1_d N_48_X1/X1/M1_g N_VDD_X1/X1/M1_s N_VDD_X1/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX2/X0/M0 N_X2/X0/6_X2/X0/M0_d N_S1_X2/X0/M0_g N_VSS_X2/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX2/X0/M1 N_16_X2/X0/M1_d N_STORE_X2/X0/M1_g N_X2/X0/6_X2/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX2/X0/M2 N_16_X2/X0/M2_d N_S1_X2/X0/M2_g N_VDD_X2/X0/M2_s N_VDD_X2/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX2/X0/M3 N_VDD_X2/X0/M3_d N_STORE_X2/X0/M3_g N_16_X2/X0/M3_s N_VDD_X2/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX2/X1/M0 N_42_X2/X1/M0_d N_16_X2/X1/M0_g N_VSS_X2/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX2/X1/M1 N_42_X2/X1/M1_d N_16_X2/X1/M1_g N_VDD_X2/X1/M1_s N_VDD_X2/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX3/X0/M0 N_X3/X0/6_X3/X0/M0_d N_19_X3/X0/M0_g N_VSS_X3/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX3/X0/M1 N_49_X3/X0/M1_d N_STATE1_X3/X0/M1_g N_X3/X0/6_X3/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX3/X0/M2 N_49_X3/X0/M2_d N_19_X3/X0/M2_g N_VDD_X3/X0/M2_s N_VDD_X3/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX3/X0/M3 N_VDD_X3/X0/M3_d N_STATE1_X3/X0/M3_g N_49_X3/X0/M3_s N_VDD_X3/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX3/X1/M0 N_MO0_X3/X1/M0_d N_49_X3/X1/M0_g N_VSS_X3/X1/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX3/X1/M1 N_MO0_X3/X1/M1_d N_49_X3/X1/M1_g N_VDD_X3/X1/M1_s N_VDD_X3/X1/M1_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX4/X0/M0 N_X4/X0/6_X4/X0/M0_d N_STATE1_X4/X0/M0_g N_VSS_X4/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX4/X0/M1 N_50_X4/X0/M1_d N_23_X4/X0/M1_g N_X4/X0/6_X4/X0/M1_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX4/X0/M2 N_50_X4/X0/M2_d N_STATE1_X4/X0/M2_g N_VDD_X4/X0/M2_s N_VDD_X4/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX4/X0/M3 N_VDD_X4/X0/M3_d N_23_X4/X0/M3_g N_50_X4/X0/M3_s N_VDD_X4/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX4/X1/M0 N_S2_X4/X1/M0_d N_50_X4/X1/M0_g N_VSS_X4/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX4/X1/M1 N_S2_X4/X1/M1_d N_50_X4/X1/M1_g N_VDD_X4/X1/M1_s N_VDD_X4/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX5/X0/M0 N_X5/X0/6_X5/X0/M0_d N_43_X5/X0/M0_g N_VSS_X5/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX5/X0/M1 N_51_X5/X0/M1_d N_POWER_X5/X0/M1_g N_X5/X0/6_X5/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX5/X0/M2 N_51_X5/X0/M2_d N_43_X5/X0/M2_g N_VDD_X5/X0/M2_s N_VDD_X5/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX5/X0/M3 N_VDD_X5/X0/M3_d N_POWER_X5/X0/M3_g N_51_X5/X0/M3_s N_VDD_X5/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX5/X1/M0 N_9_X5/X1/M0_d N_51_X5/X1/M0_g N_VSS_X5/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX5/X1/M1 N_9_X5/X1/M1_d N_51_X5/X1/M1_g N_VDD_X5/X1/M1_s N_VDD_X5/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX6/X0/M0 N_X6/X0/6_X6/X0/M0_d N_26_X6/X0/M0_g N_VSS_X6/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX6/X0/M1 N_52_X6/X0/M1_d N_STATE0_X6/X0/M1_g N_X6/X0/6_X6/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX6/X0/M2 N_52_X6/X0/M2_d N_26_X6/X0/M2_g N_VDD_X6/X0/M2_s N_VDD_X6/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX6/X0/M3 N_VDD_X6/X0/M3_d N_STATE0_X6/X0/M3_g N_52_X6/X0/M3_s N_VDD_X6/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX6/X1/M0 N_S1_X6/X1/M0_d N_52_X6/X1/M0_g N_VSS_X6/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX6/X1/M1 N_S1_X6/X1/M1_d N_52_X6/X1/M1_g N_VDD_X6/X1/M1_s N_VDD_X6/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX7/X0/M0 N_X7/X0/6_X7/X0/M0_d N_28_X7/X0/M0_g N_VSS_X7/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX7/X0/M1 N_53_X7/X0/M1_d N_STATE1_X7/X0/M1_g N_X7/X0/6_X7/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX7/X0/M2 N_53_X7/X0/M2_d N_28_X7/X0/M2_g N_VDD_X7/X0/M2_s N_VDD_X7/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX7/X0/M3 N_VDD_X7/X0/M3_d N_STATE1_X7/X0/M3_g N_53_X7/X0/M3_s N_VDD_X7/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX7/X1/M0 N_MO1_X7/X1/M0_d N_53_X7/X1/M0_g N_VSS_X7/X1/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX7/X1/M1 N_MO1_X7/X1/M1_d N_53_X7/X1/M1_g N_VDD_X7/X1/M1_s N_VDD_X7/X1/M1_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX8/X0/M0 N_X8/X0/6_X8/X0/M0_d N_16_X8/X0/M0_g N_VSS_X8/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX8/X0/M1 N_54_X8/X0/M1_d N_POWER_X8/X0/M1_g N_X8/X0/6_X8/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX8/X0/M2 N_54_X8/X0/M2_d N_16_X8/X0/M2_g N_VDD_X8/X0/M2_s N_VDD_X8/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX8/X0/M3 N_VDD_X8/X0/M3_d N_POWER_X8/X0/M3_g N_54_X8/X0/M3_s N_VDD_X8/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX8/X1/M0 N_10_X8/X1/M0_d N_54_X8/X1/M0_g N_VSS_X8/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX8/X1/M1 N_10_X8/X1/M1_d N_54_X8/X1/M1_g N_VDD_X8/X1/M1_s N_VDD_X8/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX9/X0/M0 N_X9/X0/6_X9/X0/M0_d N_26_X9/X0/M0_g N_VSS_X9/X0/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX9/X0/M1 N_55_X9/X0/M1_d N_23_X9/X0/M1_g N_X9/X0/6_X9/X0/M1_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX9/X0/M2 N_55_X9/X0/M2_d N_26_X9/X0/M2_g N_VDD_X9/X0/M2_s N_VDD_X9/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX9/X0/M3 N_VDD_X9/X0/M3_d N_23_X9/X0/M3_g N_55_X9/X0/M3_s N_VDD_X9/X0/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX9/X1/M0 N_S0_X9/X1/M0_d N_55_X9/X1/M0_g N_VSS_X9/X1/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX9/X1/M1 N_S0_X9/X1/M1_d N_55_X9/X1/M1_g N_VDD_X9/X1/M1_s N_VDD_X9/X1/M1_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX10/X0/M0 N_X10/X0/6_X10/X0/M0_d N_32_X10/X0/M0_g N_VSS_X10/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX10/X0/M1 N_56_X10/X0/M1_d N_STATE1_X10/X0/M1_g N_X10/X0/6_X10/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX10/X0/M2 N_56_X10/X0/M2_d N_32_X10/X0/M2_g N_VDD_X10/X0/M2_s N_VDD_X10/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX10/X0/M3 N_VDD_X10/X0/M3_d N_STATE1_X10/X0/M3_g N_56_X10/X0/M3_s
+ N_VDD_X10/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX10/X1/M0 N_MO2_X10/X1/M0_d N_56_X10/X1/M0_g N_VSS_X10/X1/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX10/X1/M1 N_MO2_X10/X1/M1_d N_56_X10/X1/M1_g N_VDD_X10/X1/M1_s
+ N_VDD_X10/X1/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX11/X0/M0 N_X11/X0/6_X11/X0/M0_d N_36_X11/X0/M0_g N_VSS_X11/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX11/X0/M1 N_57_X11/X0/M1_d N_STATE1_X11/X0/M1_g N_X11/X0/6_X11/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX11/X0/M2 N_57_X11/X0/M2_d N_36_X11/X0/M2_g N_VDD_X11/X0/M2_s N_VDD_X11/X0/M2_b
+ P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX11/X0/M3 N_VDD_X11/X0/M3_d N_STATE1_X11/X0/M3_g N_57_X11/X0/M3_s
+ N_VDD_X11/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX11/X1/M0 N_MO3_X11/X1/M0_d N_57_X11/X1/M0_g N_VSS_X11/X1/M0_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX11/X1/M1 N_MO3_X11/X1/M1_d N_57_X11/X1/M1_g N_VDD_X11/X1/M1_s
+ N_VDD_X11/X1/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX12/M0 N_X12/6_X12/M0_d N_42_X12/M0_g N_VSS_X12/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX12/M1 N_VSS_X12/M1_d N_S2_X12/M1_g N_X12/6_X12/M1_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX12/M2 N_X12/7_X12/M2_d N_42_X12/M2_g N_VDD_X12/M2_s N_VDD_X12/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX12/M3 N_X12/6_X12/M3_d N_S2_X12/M3_g N_X12/7_X12/M3_s N_VDD_X12/M2_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX12/X4/M0 N_43_X12/X4/M0_d N_X12/6_X12/X4/M0_g N_VSS_X12/X4/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX12/X4/M1 N_43_X12/X4/M1_d N_X12/6_X12/X4/M1_g N_VDD_X12/X4/M1_s
+ N_VDD_X12/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX13/X0/X0/M0 N_X13/X0/7_X13/X0/X0/M0_d N_12_X13/X0/X0/M0_g N_VSS_X13/X0/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX13/X0/X0/M1 N_X13/X0/7_X13/X0/X0/M1_d N_12_X13/X0/X0/M1_g N_VDD_X13/X0/X0/M1_s
+ N_VDD_X13/X0/X0/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX13/X0/X1/M0 N_X13/X0/8_X13/X0/X1/M0_d N_INIT0_X13/X0/X1/M0_g
+ N_VSS_X13/X0/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X0/X1/M1 N_X13/X0/8_X13/X0/X1/M1_d N_INIT0_X13/X0/X1/M1_g
+ N_VDD_X13/X0/X1/M1_s N_VDD_X13/X0/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X0/X2/X0/M0 N_X13/X0/X2/X0/6_X13/X0/X2/X0/M0_d N_12_X13/X0/X2/X0/M0_g
+ N_VSS_X13/X0/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX13/X0/X2/X0/M1 N_X13/X0/9_X13/X0/X2/X0/M1_d N_INIT0_X13/X0/X2/X0/M1_g
+ N_X13/X0/X2/X0/6_X13/X0/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX13/X0/X2/X0/M2 N_X13/X0/9_X13/X0/X2/X0/M2_d N_12_X13/X0/X2/X0/M2_g
+ N_VDD_X13/X0/X2/X0/M2_s N_VDD_X13/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX13/X0/X2/X0/M3 N_VDD_X13/X0/X2/X0/M3_d N_INIT0_X13/X0/X2/X0/M3_g
+ N_X13/X0/9_X13/X0/X2/X0/M3_s N_VDD_X13/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX13/X0/X2/X1/M0 N_X13/8_X13/X0/X2/X1/M0_d N_X13/X0/9_X13/X0/X2/X1/M0_g
+ N_VSS_X13/X0/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X0/X2/X1/M1 N_X13/8_X13/X0/X2/X1/M1_d N_X13/X0/9_X13/X0/X2/X1/M1_g
+ N_VDD_X13/X0/X2/X1/M1_s N_VDD_X13/X0/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X0/X3/M0 N_X13/10_X13/X0/X3/M0_d N_INIT0_X13/X0/X3/M0_g
+ N_X13/X0/7_X13/X0/X3/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X0/X3/M1 N_X13/10_X13/X0/X3/M1_d N_X13/X0/8_X13/X0/X3/M1_g
+ N_X13/X0/7_X13/X0/X3/M1_s N_VDD_X13/X0/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X0/X4/M0 N_X13/10_X13/X0/X4/M0_d N_X13/X0/8_X13/X0/X4/M0_g
+ N_12_X13/X0/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X0/X4/M1 N_X13/10_X13/X0/X4/M1_d N_INIT0_X13/X0/X4/M1_g N_12_X13/X0/X4/M1_s
+ N_VDD_X13/X0/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX13/X1/X0/M0 N_X13/X1/7_X13/X1/X0/M0_d N_X13/10_X13/X1/X0/M0_g
+ N_VSS_X13/X1/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X1/X0/M1 N_X13/X1/7_X13/X1/X0/M1_d N_X13/10_X13/X1/X0/M1_g
+ N_VDD_X13/X1/X0/M1_s N_VDD_X13/X1/X0/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X1/X1/M0 N_X13/X1/8_X13/X1/X1/M0_d N_VSS_X13/X1/X1/M0_g
+ N_VSS_X13/X1/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X1/X1/M1 N_X13/X1/8_X13/X1/X1/M1_d N_VSS_X13/X1/X1/M1_g
+ N_VDD_X13/X1/X1/M1_s N_VDD_X13/X1/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X1/X2/X0/M0 N_X13/X1/X2/X0/6_X13/X1/X2/X0/M0_d N_X13/10_X13/X1/X2/X0/M0_g
+ N_VSS_X13/X1/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX13/X1/X2/X0/M1 N_X13/X1/9_X13/X1/X2/X0/M1_d N_VSS_X13/X1/X2/X0/M1_g
+ N_X13/X1/X2/X0/6_X13/X1/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX13/X1/X2/X0/M2 N_X13/X1/9_X13/X1/X2/X0/M2_d N_X13/10_X13/X1/X2/X0/M2_g
+ N_VDD_X13/X1/X2/X0/M2_s N_VDD_X13/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX13/X1/X2/X0/M3 N_VDD_X13/X1/X2/X0/M3_d N_VSS_X13/X1/X2/X0/M3_g
+ N_X13/X1/9_X13/X1/X2/X0/M3_s N_VDD_X13/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX13/X1/X2/X1/M0 N_X13/9_X13/X1/X2/X1/M0_d N_X13/X1/9_X13/X1/X2/X1/M0_g
+ N_VSS_X13/X1/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X1/X2/X1/M1 N_X13/9_X13/X1/X2/X1/M1_d N_X13/X1/9_X13/X1/X2/X1/M1_g
+ N_VDD_X13/X1/X2/X1/M1_s N_VDD_X13/X1/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X1/X3/M0 N_2_X13/X1/X3/M0_d N_VSS_X13/X1/X3/M0_g N_X13/X1/7_X13/X1/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX13/X1/X3/M1 N_2_X13/X1/X3/M1_d N_X13/X1/8_X13/X1/X3/M1_g
+ N_X13/X1/7_X13/X1/X3/M1_s N_VDD_X13/X1/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX13/X1/X4/M0 N_2_X13/X1/X4/M0_d N_X13/X1/8_X13/X1/X4/M0_g
+ N_X13/10_X13/X1/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX13/X1/X4/M1 N_2_X13/X1/X4/M1_d N_VSS_X13/X1/X4/M1_g N_X13/10_X13/X1/X4/M1_s
+ N_VDD_X13/X1/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX13/X2/M0 N_X13/X2/6_X13/X2/M0_d N_X13/9_X13/X2/M0_g N_VSS_X13/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX13/X2/M1 N_VSS_X13/X2/M1_d N_X13/8_X13/X2/M1_g N_X13/X2/6_X13/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX13/X2/M2 N_X13/X2/7_X13/X2/M2_d N_X13/9_X13/X2/M2_g N_VDD_X13/X2/M2_s
+ N_VDD_X13/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX13/X2/M3 N_X13/X2/6_X13/X2/M3_d N_X13/8_X13/X2/M3_g N_X13/X2/7_X13/X2/M3_s
+ N_VDD_X13/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX13/X2/X4/M0 N_41_X13/X2/X4/M0_d N_X13/X2/6_X13/X2/X4/M0_g N_VSS_X13/X2/X4/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX13/X2/X4/M1 N_41_X13/X2/X4/M1_d N_X13/X2/6_X13/X2/X4/M1_g N_VDD_X13/X2/X4/M1_s
+ N_VDD_X13/X2/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX14/X0/X0/M0 N_X14/X0/7_X14/X0/X0/M0_d N_24_X14/X0/X0/M0_g N_VSS_X14/X0/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX14/X0/X0/M1 N_X14/X0/7_X14/X0/X0/M1_d N_24_X14/X0/X0/M1_g N_VDD_X14/X0/X0/M1_s
+ N_VDD_X14/X0/X0/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX14/X0/X1/M0 N_X14/X0/8_X14/X0/X1/M0_d N_INIT1_X14/X0/X1/M0_g
+ N_VSS_X14/X0/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X0/X1/M1 N_X14/X0/8_X14/X0/X1/M1_d N_INIT1_X14/X0/X1/M1_g
+ N_VDD_X14/X0/X1/M1_s N_VDD_X14/X0/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X0/X2/X0/M0 N_X14/X0/X2/X0/6_X14/X0/X2/X0/M0_d N_24_X14/X0/X2/X0/M0_g
+ N_VSS_X14/X0/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX14/X0/X2/X0/M1 N_X14/X0/9_X14/X0/X2/X0/M1_d N_INIT1_X14/X0/X2/X0/M1_g
+ N_X14/X0/X2/X0/6_X14/X0/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX14/X0/X2/X0/M2 N_X14/X0/9_X14/X0/X2/X0/M2_d N_24_X14/X0/X2/X0/M2_g
+ N_VDD_X14/X0/X2/X0/M2_s N_VDD_X14/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX14/X0/X2/X0/M3 N_VDD_X14/X0/X2/X0/M3_d N_INIT1_X14/X0/X2/X0/M3_g
+ N_X14/X0/9_X14/X0/X2/X0/M3_s N_VDD_X14/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX14/X0/X2/X1/M0 N_X14/8_X14/X0/X2/X1/M0_d N_X14/X0/9_X14/X0/X2/X1/M0_g
+ N_VSS_X14/X0/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X0/X2/X1/M1 N_X14/8_X14/X0/X2/X1/M1_d N_X14/X0/9_X14/X0/X2/X1/M1_g
+ N_VDD_X14/X0/X2/X1/M1_s N_VDD_X14/X0/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X0/X3/M0 N_X14/10_X14/X0/X3/M0_d N_INIT1_X14/X0/X3/M0_g
+ N_X14/X0/7_X14/X0/X3/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X0/X3/M1 N_X14/10_X14/X0/X3/M1_d N_X14/X0/8_X14/X0/X3/M1_g
+ N_X14/X0/7_X14/X0/X3/M1_s N_VDD_X14/X0/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X0/X4/M0 N_X14/10_X14/X0/X4/M0_d N_X14/X0/8_X14/X0/X4/M0_g
+ N_24_X14/X0/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X0/X4/M1 N_X14/10_X14/X0/X4/M1_d N_INIT1_X14/X0/X4/M1_g N_24_X14/X0/X4/M1_s
+ N_VDD_X14/X0/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX14/X1/X0/M0 N_X14/X1/7_X14/X1/X0/M0_d N_X14/10_X14/X1/X0/M0_g
+ N_VSS_X14/X1/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X1/X0/M1 N_X14/X1/7_X14/X1/X0/M1_d N_X14/10_X14/X1/X0/M1_g
+ N_VDD_X14/X1/X0/M1_s N_VDD_X14/X1/X0/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X1/X1/M0 N_X14/X1/8_X14/X1/X1/M0_d N_41_X14/X1/X1/M0_g N_VSS_X14/X1/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX14/X1/X1/M1 N_X14/X1/8_X14/X1/X1/M1_d N_41_X14/X1/X1/M1_g N_VDD_X14/X1/X1/M1_s
+ N_VDD_X14/X1/X1/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX14/X1/X2/X0/M0 N_X14/X1/X2/X0/6_X14/X1/X2/X0/M0_d N_X14/10_X14/X1/X2/X0/M0_g
+ N_VSS_X14/X1/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX14/X1/X2/X0/M1 N_X14/X1/9_X14/X1/X2/X0/M1_d N_41_X14/X1/X2/X0/M1_g
+ N_X14/X1/X2/X0/6_X14/X1/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX14/X1/X2/X0/M2 N_X14/X1/9_X14/X1/X2/X0/M2_d N_X14/10_X14/X1/X2/X0/M2_g
+ N_VDD_X14/X1/X2/X0/M2_s N_VDD_X14/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX14/X1/X2/X0/M3 N_VDD_X14/X1/X2/X0/M3_d N_41_X14/X1/X2/X0/M3_g
+ N_X14/X1/9_X14/X1/X2/X0/M3_s N_VDD_X14/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX14/X1/X2/X1/M0 N_X14/9_X14/X1/X2/X1/M0_d N_X14/X1/9_X14/X1/X2/X1/M0_g
+ N_VSS_X14/X1/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X1/X2/X1/M1 N_X14/9_X14/X1/X2/X1/M1_d N_X14/X1/9_X14/X1/X2/X1/M1_g
+ N_VDD_X14/X1/X2/X1/M1_s N_VDD_X14/X1/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X1/X3/M0 N_4_X14/X1/X3/M0_d N_41_X14/X1/X3/M0_g N_X14/X1/7_X14/X1/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX14/X1/X3/M1 N_4_X14/X1/X3/M1_d N_X14/X1/8_X14/X1/X3/M1_g
+ N_X14/X1/7_X14/X1/X3/M1_s N_VDD_X14/X1/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX14/X1/X4/M0 N_4_X14/X1/X4/M0_d N_X14/X1/8_X14/X1/X4/M0_g
+ N_X14/10_X14/X1/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX14/X1/X4/M1 N_4_X14/X1/X4/M1_d N_41_X14/X1/X4/M1_g N_X14/10_X14/X1/X4/M1_s
+ N_VDD_X14/X1/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX14/X2/M0 N_X14/X2/6_X14/X2/M0_d N_X14/9_X14/X2/M0_g N_VSS_X14/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX14/X2/M1 N_VSS_X14/X2/M1_d N_X14/8_X14/X2/M1_g N_X14/X2/6_X14/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX14/X2/M2 N_X14/X2/7_X14/X2/M2_d N_X14/9_X14/X2/M2_g N_VDD_X14/X2/M2_s
+ N_VDD_X14/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX14/X2/M3 N_X14/X2/6_X14/X2/M3_d N_X14/8_X14/X2/M3_g N_X14/X2/7_X14/X2/M3_s
+ N_VDD_X14/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX14/X2/X4/M0 N_44_X14/X2/X4/M0_d N_X14/X2/6_X14/X2/X4/M0_g N_VSS_X14/X2/X4/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX14/X2/X4/M1 N_44_X14/X2/X4/M1_d N_X14/X2/6_X14/X2/X4/M1_g N_VDD_X14/X2/X4/M1_s
+ N_VDD_X14/X2/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX15/X0/X0/M0 N_X15/X0/7_X15/X0/X0/M0_d N_31_X15/X0/X0/M0_g N_VSS_X15/X0/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX15/X0/X0/M1 N_X15/X0/7_X15/X0/X0/M1_d N_31_X15/X0/X0/M1_g N_VDD_X15/X0/X0/M1_s
+ N_VDD_X15/X0/X0/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX15/X0/X1/M0 N_X15/X0/8_X15/X0/X1/M0_d N_INIT2_X15/X0/X1/M0_g
+ N_VSS_X15/X0/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X0/X1/M1 N_X15/X0/8_X15/X0/X1/M1_d N_INIT2_X15/X0/X1/M1_g
+ N_VDD_X15/X0/X1/M1_s N_VDD_X15/X0/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X0/X2/X0/M0 N_X15/X0/X2/X0/6_X15/X0/X2/X0/M0_d N_31_X15/X0/X2/X0/M0_g
+ N_VSS_X15/X0/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX15/X0/X2/X0/M1 N_X15/X0/9_X15/X0/X2/X0/M1_d N_INIT2_X15/X0/X2/X0/M1_g
+ N_X15/X0/X2/X0/6_X15/X0/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX15/X0/X2/X0/M2 N_X15/X0/9_X15/X0/X2/X0/M2_d N_31_X15/X0/X2/X0/M2_g
+ N_VDD_X15/X0/X2/X0/M2_s N_VDD_X15/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX15/X0/X2/X0/M3 N_VDD_X15/X0/X2/X0/M3_d N_INIT2_X15/X0/X2/X0/M3_g
+ N_X15/X0/9_X15/X0/X2/X0/M3_s N_VDD_X15/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX15/X0/X2/X1/M0 N_X15/8_X15/X0/X2/X1/M0_d N_X15/X0/9_X15/X0/X2/X1/M0_g
+ N_VSS_X15/X0/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X0/X2/X1/M1 N_X15/8_X15/X0/X2/X1/M1_d N_X15/X0/9_X15/X0/X2/X1/M1_g
+ N_VDD_X15/X0/X2/X1/M1_s N_VDD_X15/X0/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X0/X3/M0 N_X15/10_X15/X0/X3/M0_d N_INIT2_X15/X0/X3/M0_g
+ N_X15/X0/7_X15/X0/X3/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X0/X3/M1 N_X15/10_X15/X0/X3/M1_d N_X15/X0/8_X15/X0/X3/M1_g
+ N_X15/X0/7_X15/X0/X3/M1_s N_VDD_X15/X0/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X0/X4/M0 N_X15/10_X15/X0/X4/M0_d N_X15/X0/8_X15/X0/X4/M0_g
+ N_31_X15/X0/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X0/X4/M1 N_X15/10_X15/X0/X4/M1_d N_INIT2_X15/X0/X4/M1_g N_31_X15/X0/X4/M1_s
+ N_VDD_X15/X0/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX15/X1/X0/M0 N_X15/X1/7_X15/X1/X0/M0_d N_X15/10_X15/X1/X0/M0_g
+ N_VSS_X15/X1/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X1/X0/M1 N_X15/X1/7_X15/X1/X0/M1_d N_X15/10_X15/X1/X0/M1_g
+ N_VDD_X15/X1/X0/M1_s N_VDD_X15/X1/X0/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X1/X1/M0 N_X15/X1/8_X15/X1/X1/M0_d N_44_X15/X1/X1/M0_g N_VSS_X15/X1/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX15/X1/X1/M1 N_X15/X1/8_X15/X1/X1/M1_d N_44_X15/X1/X1/M1_g N_VDD_X15/X1/X1/M1_s
+ N_VDD_X15/X1/X1/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX15/X1/X2/X0/M0 N_X15/X1/X2/X0/6_X15/X1/X2/X0/M0_d N_X15/10_X15/X1/X2/X0/M0_g
+ N_VSS_X15/X1/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX15/X1/X2/X0/M1 N_X15/X1/9_X15/X1/X2/X0/M1_d N_44_X15/X1/X2/X0/M1_g
+ N_X15/X1/X2/X0/6_X15/X1/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX15/X1/X2/X0/M2 N_X15/X1/9_X15/X1/X2/X0/M2_d N_X15/10_X15/X1/X2/X0/M2_g
+ N_VDD_X15/X1/X2/X0/M2_s N_VDD_X15/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX15/X1/X2/X0/M3 N_VDD_X15/X1/X2/X0/M3_d N_44_X15/X1/X2/X0/M3_g
+ N_X15/X1/9_X15/X1/X2/X0/M3_s N_VDD_X15/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX15/X1/X2/X1/M0 N_X15/9_X15/X1/X2/X1/M0_d N_X15/X1/9_X15/X1/X2/X1/M0_g
+ N_VSS_X15/X1/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X1/X2/X1/M1 N_X15/9_X15/X1/X2/X1/M1_d N_X15/X1/9_X15/X1/X2/X1/M1_g
+ N_VDD_X15/X1/X2/X1/M1_s N_VDD_X15/X1/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X1/X3/M0 N_6_X15/X1/X3/M0_d N_44_X15/X1/X3/M0_g N_X15/X1/7_X15/X1/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX15/X1/X3/M1 N_6_X15/X1/X3/M1_d N_X15/X1/8_X15/X1/X3/M1_g
+ N_X15/X1/7_X15/X1/X3/M1_s N_VDD_X15/X1/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX15/X1/X4/M0 N_6_X15/X1/X4/M0_d N_X15/X1/8_X15/X1/X4/M0_g
+ N_X15/10_X15/X1/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX15/X1/X4/M1 N_6_X15/X1/X4/M1_d N_44_X15/X1/X4/M1_g N_X15/10_X15/X1/X4/M1_s
+ N_VDD_X15/X1/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX15/X2/M0 N_X15/X2/6_X15/X2/M0_d N_X15/9_X15/X2/M0_g N_VSS_X15/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX15/X2/M1 N_VSS_X15/X2/M1_d N_X15/8_X15/X2/M1_g N_X15/X2/6_X15/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX15/X2/M2 N_X15/X2/7_X15/X2/M2_d N_X15/9_X15/X2/M2_g N_VDD_X15/X2/M2_s
+ N_VDD_X15/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX15/X2/M3 N_X15/X2/6_X15/X2/M3_d N_X15/8_X15/X2/M3_g N_X15/X2/7_X15/X2/M3_s
+ N_VDD_X15/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX15/X2/X4/M0 N_46_X15/X2/X4/M0_d N_X15/X2/6_X15/X2/X4/M0_g N_VSS_X15/X2/X4/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX15/X2/X4/M1 N_46_X15/X2/X4/M1_d N_X15/X2/6_X15/X2/X4/M1_g N_VDD_X15/X2/X4/M1_s
+ N_VDD_X15/X2/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX16/X0/X0/M0 N_X16/X0/7_X16/X0/X0/M0_d N_35_X16/X0/X0/M0_g N_VSS_X16/X0/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX16/X0/X0/M1 N_X16/X0/7_X16/X0/X0/M1_d N_35_X16/X0/X0/M1_g N_VDD_X16/X0/X0/M1_s
+ N_VDD_X16/X0/X0/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX16/X0/X1/M0 N_X16/X0/8_X16/X0/X1/M0_d N_INIT3_X16/X0/X1/M0_g
+ N_VSS_X16/X0/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X0/X1/M1 N_X16/X0/8_X16/X0/X1/M1_d N_INIT3_X16/X0/X1/M1_g
+ N_VDD_X16/X0/X1/M1_s N_VDD_X16/X0/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X0/X2/X0/M0 N_X16/X0/X2/X0/6_X16/X0/X2/X0/M0_d N_35_X16/X0/X2/X0/M0_g
+ N_VSS_X16/X0/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX16/X0/X2/X0/M1 N_X16/X0/9_X16/X0/X2/X0/M1_d N_INIT3_X16/X0/X2/X0/M1_g
+ N_X16/X0/X2/X0/6_X16/X0/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX16/X0/X2/X0/M2 N_X16/X0/9_X16/X0/X2/X0/M2_d N_35_X16/X0/X2/X0/M2_g
+ N_VDD_X16/X0/X2/X0/M2_s N_VDD_X16/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX16/X0/X2/X0/M3 N_VDD_X16/X0/X2/X0/M3_d N_INIT3_X16/X0/X2/X0/M3_g
+ N_X16/X0/9_X16/X0/X2/X0/M3_s N_VDD_X16/X0/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX16/X0/X2/X1/M0 N_X16/8_X16/X0/X2/X1/M0_d N_X16/X0/9_X16/X0/X2/X1/M0_g
+ N_VSS_X16/X0/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X0/X2/X1/M1 N_X16/8_X16/X0/X2/X1/M1_d N_X16/X0/9_X16/X0/X2/X1/M1_g
+ N_VDD_X16/X0/X2/X1/M1_s N_VDD_X16/X0/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X0/X3/M0 N_X16/10_X16/X0/X3/M0_d N_INIT3_X16/X0/X3/M0_g
+ N_X16/X0/7_X16/X0/X3/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X0/X3/M1 N_X16/10_X16/X0/X3/M1_d N_X16/X0/8_X16/X0/X3/M1_g
+ N_X16/X0/7_X16/X0/X3/M1_s N_VDD_X16/X0/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X0/X4/M0 N_X16/10_X16/X0/X4/M0_d N_X16/X0/8_X16/X0/X4/M0_g
+ N_35_X16/X0/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X0/X4/M1 N_X16/10_X16/X0/X4/M1_d N_INIT3_X16/X0/X4/M1_g N_35_X16/X0/X4/M1_s
+ N_VDD_X16/X0/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX16/X1/X0/M0 N_X16/X1/7_X16/X1/X0/M0_d N_X16/10_X16/X1/X0/M0_g
+ N_VSS_X16/X1/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X1/X0/M1 N_X16/X1/7_X16/X1/X0/M1_d N_X16/10_X16/X1/X0/M1_g
+ N_VDD_X16/X1/X0/M1_s N_VDD_X16/X1/X0/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X1/X1/M0 N_X16/X1/8_X16/X1/X1/M0_d N_46_X16/X1/X1/M0_g N_VSS_X16/X1/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX16/X1/X1/M1 N_X16/X1/8_X16/X1/X1/M1_d N_46_X16/X1/X1/M1_g N_VDD_X16/X1/X1/M1_s
+ N_VDD_X16/X1/X1/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX16/X1/X2/X0/M0 N_X16/X1/X2/X0/6_X16/X1/X2/X0/M0_d N_X16/10_X16/X1/X2/X0/M0_g
+ N_VSS_X16/X1/X2/X0/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX16/X1/X2/X0/M1 N_X16/X1/9_X16/X1/X2/X0/M1_d N_46_X16/X1/X2/X0/M1_g
+ N_X16/X1/X2/X0/6_X16/X1/X2/X0/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX16/X1/X2/X0/M2 N_X16/X1/9_X16/X1/X2/X0/M2_d N_X16/10_X16/X1/X2/X0/M2_g
+ N_VDD_X16/X1/X2/X0/M2_s N_VDD_X16/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX16/X1/X2/X0/M3 N_VDD_X16/X1/X2/X0/M3_d N_46_X16/X1/X2/X0/M3_g
+ N_X16/X1/9_X16/X1/X2/X0/M3_s N_VDD_X16/X1/X2/X0/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX16/X1/X2/X1/M0 N_X16/9_X16/X1/X2/X1/M0_d N_X16/X1/9_X16/X1/X2/X1/M0_g
+ N_VSS_X16/X1/X2/X1/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X1/X2/X1/M1 N_X16/9_X16/X1/X2/X1/M1_d N_X16/X1/9_X16/X1/X2/X1/M1_g
+ N_VDD_X16/X1/X2/X1/M1_s N_VDD_X16/X1/X2/X1/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X1/X3/M0 N_8_X16/X1/X3/M0_d N_46_X16/X1/X3/M0_g N_X16/X1/7_X16/X1/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX16/X1/X3/M1 N_8_X16/X1/X3/M1_d N_X16/X1/8_X16/X1/X3/M1_g
+ N_X16/X1/7_X16/X1/X3/M1_s N_VDD_X16/X1/X3/M1_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=2.275e-12 PD=4.32e-06 PS=4.32e-06
mX16/X1/X4/M0 N_8_X16/X1/X4/M0_d N_X16/X1/8_X16/X1/X4/M0_g
+ N_X16/10_X16/X1/X4/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13
+ AS=9.1e-13 PD=2.82e-06 PS=2.82e-06
mX16/X1/X4/M1 N_8_X16/X1/X4/M1_d N_46_X16/X1/X4/M1_g N_X16/10_X16/X1/X4/M1_s
+ N_VDD_X16/X1/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX16/X2/M0 N_X16/X2/6_X16/X2/M0_d N_X16/9_X16/X2/M0_g N_VSS_X16/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX16/X2/M1 N_VSS_X16/X2/M1_d N_X16/8_X16/X2/M1_g N_X16/X2/6_X16/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX16/X2/M2 N_X16/X2/7_X16/X2/M2_d N_X16/9_X16/X2/M2_g N_VDD_X16/X2/M2_s
+ N_VDD_X16/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX16/X2/M3 N_X16/X2/6_X16/X2/M3_d N_X16/8_X16/X2/M3_g N_X16/X2/7_X16/X2/M3_s
+ N_VDD_X16/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX16/X2/X4/M0 N_58_X16/X2/X4/M0_d N_X16/X2/6_X16/X2/X4/M0_g N_VSS_X16/X2/X4/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX16/X2/X4/M1 N_58_X16/X2/X4/M1_d N_X16/X2/6_X16/X2/X4/M1_g N_VDD_X16/X2/X4/M1_s
+ N_VDD_X16/X2/X4/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX17/M0 N_X17/11_X17/M0_d N_X17/7_X17/M0_g N_VSS_X17/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX17/M1 N_X17/12_X17/M1_d N_CLK_X17/M1_g N_X17/11_X17/M1_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07 PS=8.2e-07
mX17/M2 N_X17/9_X17/M2_d N_X17/8_X17/M2_g N_X17/12_X17/M2_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX17/M3 N_X17/9_X17/M3_d N_X17/7_X17/M3_g N_VDD_X17/M3_s N_VDD_X17/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX17/M4 N_VDD_X17/M4_d N_CLK_X17/M4_g N_X17/9_X17/M4_s N_VDD_X17/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12 PD=8.2e-07 PS=8.2e-07
mX17/M5 N_X17/9_X17/M5_d N_X17/8_X17/M5_g N_VDD_X17/M5_s N_VDD_X17/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX17/X6/M0 N_X17/X6/6_X17/X6/M0_d N_X17/8_X17/X6/M0_g N_VSS_X17/X6/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX17/X6/M1 N_X17/10_X17/X6/M1_d N_X17/7_X17/X6/M1_g N_X17/X6/6_X17/X6/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX17/X6/M2 N_X17/10_X17/X6/M2_d N_X17/8_X17/X6/M2_g N_VDD_X17/X6/M2_s
+ N_VDD_X17/X6/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX17/X6/M3 N_VDD_X17/X6/M3_d N_X17/7_X17/X6/M3_g N_X17/10_X17/X6/M3_s
+ N_VDD_X17/X6/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX17/X7/M0 N_X17/X7/6_X17/X7/M0_d N_X17/10_X17/X7/M0_g N_VSS_X17/X7/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX17/X7/M1 N_X17/7_X17/X7/M1_d N_CLK_X17/X7/M1_g N_X17/X7/6_X17/X7/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX17/X7/M2 N_X17/7_X17/X7/M2_d N_X17/10_X17/X7/M2_g N_VDD_X17/X7/M2_s
+ N_VDD_X17/X7/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX17/X7/M3 N_VDD_X17/X7/M3_d N_CLK_X17/X7/M3_g N_X17/7_X17/X7/M3_s
+ N_VDD_X17/X7/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX17/X8/M0 N_X17/X8/6_X17/X8/M0_d N_X17/7_X17/X8/M0_g N_VSS_X17/X8/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX17/X8/M1 N_STATE0_X17/X8/M1_d N_23_X17/X8/M1_g N_X17/X8/6_X17/X8/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX17/X8/M2 N_STATE0_X17/X8/M2_d N_X17/7_X17/X8/M2_g N_VDD_X17/X8/M2_s
+ N_VDD_X17/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX17/X8/M3 N_VDD_X17/X8/M3_d N_23_X17/X8/M3_g N_STATE0_X17/X8/M3_s
+ N_VDD_X17/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX17/X9/M0 N_X17/X9/6_X17/X9/M0_d N_STATE0_X17/X9/M0_g N_VSS_X17/X9/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX17/X9/M1 N_23_X17/X9/M1_d N_X17/9_X17/X9/M1_g N_X17/X9/6_X17/X9/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX17/X9/M2 N_23_X17/X9/M2_d N_STATE0_X17/X9/M2_g N_VDD_X17/X9/M2_s
+ N_VDD_X17/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX17/X9/M3 N_VDD_X17/X9/M3_d N_X17/9_X17/X9/M3_g N_23_X17/X9/M3_s
+ N_VDD_X17/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX17/X10/M0 N_X17/X10/6_X17/X10/M0_d N_X17/9_X17/X10/M0_g N_VSS_X17/X10/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX17/X10/M1 N_X17/8_X17/X10/M1_d N_10_X17/X10/M1_g N_X17/X10/6_X17/X10/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX17/X10/M2 N_X17/8_X17/X10/M2_d N_X17/9_X17/X10/M2_g N_VDD_X17/X10/M2_s
+ N_VDD_X17/X10/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX17/X10/M3 N_VDD_X17/X10/M3_d N_10_X17/X10/M3_g N_X17/8_X17/X10/M3_s
+ N_VDD_X17/X10/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX18/M0 N_X18/11_X18/M0_d N_X18/7_X18/M0_g N_VSS_X18/M0_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX18/M1 N_X18/12_X18/M1_d N_CLK_X18/M1_g N_X18/11_X18/M1_s N_VSS_X0/X0/M0_b N_18
+ L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07 PS=8.2e-07
mX18/M2 N_X18/9_X18/M2_d N_X18/8_X18/M2_g N_X18/12_X18/M2_s N_VSS_X0/X0/M0_b
+ N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX18/M3 N_X18/9_X18/M3_d N_X18/7_X18/M3_g N_VDD_X18/M3_s N_VDD_X18/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX18/M4 N_VDD_X18/M4_d N_CLK_X18/M4_g N_X18/9_X18/M4_s N_VDD_X18/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12 PD=8.2e-07 PS=8.2e-07
mX18/M5 N_X18/9_X18/M5_d N_X18/8_X18/M5_g N_VDD_X18/M5_s N_VDD_X18/M3_b P_18
+ L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX18/X6/M0 N_X18/X6/6_X18/X6/M0_d N_X18/8_X18/X6/M0_g N_VSS_X18/X6/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX18/X6/M1 N_X18/10_X18/X6/M1_d N_X18/7_X18/X6/M1_g N_X18/X6/6_X18/X6/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX18/X6/M2 N_X18/10_X18/X6/M2_d N_X18/8_X18/X6/M2_g N_VDD_X18/X6/M2_s
+ N_VDD_X18/X6/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX18/X6/M3 N_VDD_X18/X6/M3_d N_X18/7_X18/X6/M3_g N_X18/10_X18/X6/M3_s
+ N_VDD_X18/X6/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX18/X7/M0 N_X18/X7/6_X18/X7/M0_d N_X18/10_X18/X7/M0_g N_VSS_X18/X7/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX18/X7/M1 N_X18/7_X18/X7/M1_d N_CLK_X18/X7/M1_g N_X18/X7/6_X18/X7/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX18/X7/M2 N_X18/7_X18/X7/M2_d N_X18/10_X18/X7/M2_g N_VDD_X18/X7/M2_s
+ N_VDD_X18/X7/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX18/X7/M3 N_VDD_X18/X7/M3_d N_CLK_X18/X7/M3_g N_X18/7_X18/X7/M3_s
+ N_VDD_X18/X7/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX18/X8/M0 N_X18/X8/6_X18/X8/M0_d N_X18/7_X18/X8/M0_g N_VSS_X18/X8/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX18/X8/M1 N_STATE1_X18/X8/M1_d N_26_X18/X8/M1_g N_X18/X8/6_X18/X8/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX18/X8/M2 N_STATE1_X18/X8/M2_d N_X18/7_X18/X8/M2_g N_VDD_X18/X8/M2_s
+ N_VDD_X18/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX18/X8/M3 N_VDD_X18/X8/M3_d N_26_X18/X8/M3_g N_STATE1_X18/X8/M3_s
+ N_VDD_X18/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX18/X9/M0 N_X18/X9/6_X18/X9/M0_d N_STATE1_X18/X9/M0_g N_VSS_X18/X9/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX18/X9/M1 N_26_X18/X9/M1_d N_X18/9_X18/X9/M1_g N_X18/X9/6_X18/X9/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX18/X9/M2 N_26_X18/X9/M2_d N_STATE1_X18/X9/M2_g N_VDD_X18/X9/M2_s
+ N_VDD_X18/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX18/X9/M3 N_VDD_X18/X9/M3_d N_X18/9_X18/X9/M3_g N_26_X18/X9/M3_s
+ N_VDD_X18/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX18/X10/M0 N_X18/X10/6_X18/X10/M0_d N_X18/9_X18/X10/M0_g N_VSS_X18/X10/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX18/X10/M1 N_X18/8_X18/X10/M1_d N_9_X18/X10/M1_g N_X18/X10/6_X18/X10/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX18/X10/M2 N_X18/8_X18/X10/M2_d N_X18/9_X18/X10/M2_g N_VDD_X18/X10/M2_s
+ N_VDD_X18/X10/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX18/X10/M3 N_VDD_X18/X10/M3_d N_9_X18/X10/M3_g N_X18/8_X18/X10/M3_s
+ N_VDD_X18/X10/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX19/X0/M0 N_X19/X0/6_X19/X0/M0_d N_X19/8_X19/X0/M0_g N_VSS_X19/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX19/X0/M1 N_X19/7_X19/X0/M1_d N_INIT0_X19/X0/M1_g N_X19/X0/6_X19/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX19/X0/M2 N_X19/7_X19/X0/M2_d N_X19/8_X19/X0/M2_g N_VDD_X19/X0/M2_s
+ N_VDD_X19/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX19/X0/M3 N_VDD_X19/X0/M3_d N_INIT0_X19/X0/M3_g N_X19/7_X19/X0/M3_s
+ N_VDD_X19/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX19/X1/M0 N_X19/X1/6_X19/X1/M0_d N_11_X19/X1/M0_g N_VSS_X19/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX19/X1/M1 N_X19/9_X19/X1/M1_d N_2_X19/X1/M1_g N_X19/X1/6_X19/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX19/X1/M2 N_X19/9_X19/X1/M2_d N_11_X19/X1/M2_g N_VDD_X19/X1/M2_s
+ N_VDD_X19/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX19/X1/M3 N_VDD_X19/X1/M3_d N_2_X19/X1/M3_g N_X19/9_X19/X1/M3_s
+ N_VDD_X19/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX19/X2/M0 N_X19/X2/6_X19/X2/M0_d N_X19/9_X19/X2/M0_g N_VSS_X19/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX19/X2/M1 N_17_X19/X2/M1_d N_X19/7_X19/X2/M1_g N_X19/X2/6_X19/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX19/X2/M2 N_17_X19/X2/M2_d N_X19/9_X19/X2/M2_g N_VDD_X19/X2/M2_s
+ N_VDD_X19/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX19/X2/M3 N_VDD_X19/X2/M3_d N_X19/7_X19/X2/M3_g N_17_X19/X2/M3_s
+ N_VDD_X19/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX19/X3/M0 N_X19/8_X19/X3/M0_d N_11_X19/X3/M0_g N_VSS_X19/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX19/X3/M1 N_X19/8_X19/X3/M1_d N_11_X19/X3/M1_g N_VDD_X19/X3/M1_s
+ N_VDD_X19/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX20/X0/M0 N_X20/X0/6_X20/X0/M0_d N_X20/8_X20/X0/M0_g N_VSS_X20/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX20/X0/M1 N_X20/7_X20/X0/M1_d N_12_X20/X0/M1_g N_X20/X0/6_X20/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX20/X0/M2 N_X20/7_X20/X0/M2_d N_X20/8_X20/X0/M2_g N_VDD_X20/X0/M2_s
+ N_VDD_X20/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX20/X0/M3 N_VDD_X20/X0/M3_d N_12_X20/X0/M3_g N_X20/7_X20/X0/M3_s
+ N_VDD_X20/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX20/X1/M0 N_X20/X1/6_X20/X1/M0_d N_STATE0_X20/X1/M0_g N_VSS_X20/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX20/X1/M1 N_X20/9_X20/X1/M1_d N_INIT0_X20/X1/M1_g N_X20/X1/6_X20/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX20/X1/M2 N_X20/9_X20/X1/M2_d N_STATE0_X20/X1/M2_g N_VDD_X20/X1/M2_s
+ N_VDD_X20/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX20/X1/M3 N_VDD_X20/X1/M3_d N_INIT0_X20/X1/M3_g N_X20/9_X20/X1/M3_s
+ N_VDD_X20/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX20/X2/M0 N_X20/X2/6_X20/X2/M0_d N_X20/9_X20/X2/M0_g N_VSS_X20/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX20/X2/M1 N_19_X20/X2/M1_d N_X20/7_X20/X2/M1_g N_X20/X2/6_X20/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX20/X2/M2 N_19_X20/X2/M2_d N_X20/9_X20/X2/M2_g N_VDD_X20/X2/M2_s
+ N_VDD_X20/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX20/X2/M3 N_VDD_X20/X2/M3_d N_X20/7_X20/X2/M3_g N_19_X20/X2/M3_s
+ N_VDD_X20/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX20/X3/M0 N_X20/8_X20/X3/M0_d N_STATE0_X20/X3/M0_g N_VSS_X20/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX20/X3/M1 N_X20/8_X20/X3/M1_d N_STATE0_X20/X3/M1_g N_VDD_X20/X3/M1_s
+ N_VDD_X20/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX21/X0/M0 N_X21/X0/6_X21/X0/M0_d N_X21/8_X21/X0/M0_g N_VSS_X21/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX21/X0/M1 N_X21/7_X21/X0/M1_d N_INIT1_X21/X0/M1_g N_X21/X0/6_X21/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX21/X0/M2 N_X21/7_X21/X0/M2_d N_X21/8_X21/X0/M2_g N_VDD_X21/X0/M2_s
+ N_VDD_X21/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX21/X0/M3 N_VDD_X21/X0/M3_d N_INIT1_X21/X0/M3_g N_X21/7_X21/X0/M3_s
+ N_VDD_X21/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX21/X1/M0 N_X21/X1/6_X21/X1/M0_d N_11_X21/X1/M0_g N_VSS_X21/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX21/X1/M1 N_X21/9_X21/X1/M1_d N_4_X21/X1/M1_g N_X21/X1/6_X21/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX21/X1/M2 N_X21/9_X21/X1/M2_d N_11_X21/X1/M2_g N_VDD_X21/X1/M2_s
+ N_VDD_X21/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX21/X1/M3 N_VDD_X21/X1/M3_d N_4_X21/X1/M3_g N_X21/9_X21/X1/M3_s
+ N_VDD_X21/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX21/X2/M0 N_X21/X2/6_X21/X2/M0_d N_X21/9_X21/X2/M0_g N_VSS_X21/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX21/X2/M1 N_27_X21/X2/M1_d N_X21/7_X21/X2/M1_g N_X21/X2/6_X21/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX21/X2/M2 N_27_X21/X2/M2_d N_X21/9_X21/X2/M2_g N_VDD_X21/X2/M2_s
+ N_VDD_X21/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX21/X2/M3 N_VDD_X21/X2/M3_d N_X21/7_X21/X2/M3_g N_27_X21/X2/M3_s
+ N_VDD_X21/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX21/X3/M0 N_X21/8_X21/X3/M0_d N_11_X21/X3/M0_g N_VSS_X21/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX21/X3/M1 N_X21/8_X21/X3/M1_d N_11_X21/X3/M1_g N_VDD_X21/X3/M1_s
+ N_VDD_X21/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX22/X0/M0 N_X22/X0/6_X22/X0/M0_d N_X22/8_X22/X0/M0_g N_VSS_X22/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX22/X0/M1 N_X22/7_X22/X0/M1_d N_24_X22/X0/M1_g N_X22/X0/6_X22/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX22/X0/M2 N_X22/7_X22/X0/M2_d N_X22/8_X22/X0/M2_g N_VDD_X22/X0/M2_s
+ N_VDD_X22/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX22/X0/M3 N_VDD_X22/X0/M3_d N_24_X22/X0/M3_g N_X22/7_X22/X0/M3_s
+ N_VDD_X22/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX22/X1/M0 N_X22/X1/6_X22/X1/M0_d N_STATE0_X22/X1/M0_g N_VSS_X22/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX22/X1/M1 N_X22/9_X22/X1/M1_d N_INIT1_X22/X1/M1_g N_X22/X1/6_X22/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX22/X1/M2 N_X22/9_X22/X1/M2_d N_STATE0_X22/X1/M2_g N_VDD_X22/X1/M2_s
+ N_VDD_X22/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX22/X1/M3 N_VDD_X22/X1/M3_d N_INIT1_X22/X1/M3_g N_X22/9_X22/X1/M3_s
+ N_VDD_X22/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX22/X2/M0 N_X22/X2/6_X22/X2/M0_d N_X22/9_X22/X2/M0_g N_VSS_X22/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX22/X2/M1 N_28_X22/X2/M1_d N_X22/7_X22/X2/M1_g N_X22/X2/6_X22/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX22/X2/M2 N_28_X22/X2/M2_d N_X22/9_X22/X2/M2_g N_VDD_X22/X2/M2_s
+ N_VDD_X22/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX22/X2/M3 N_VDD_X22/X2/M3_d N_X22/7_X22/X2/M3_g N_28_X22/X2/M3_s
+ N_VDD_X22/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX22/X3/M0 N_X22/8_X22/X3/M0_d N_STATE0_X22/X3/M0_g N_VSS_X22/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX22/X3/M1 N_X22/8_X22/X3/M1_d N_STATE0_X22/X3/M1_g N_VDD_X22/X3/M1_s
+ N_VDD_X22/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX23/X0/M0 N_X23/X0/6_X23/X0/M0_d N_X23/8_X23/X0/M0_g N_VSS_X23/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX23/X0/M1 N_X23/7_X23/X0/M1_d N_31_X23/X0/M1_g N_X23/X0/6_X23/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX23/X0/M2 N_X23/7_X23/X0/M2_d N_X23/8_X23/X0/M2_g N_VDD_X23/X0/M2_s
+ N_VDD_X23/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX23/X0/M3 N_VDD_X23/X0/M3_d N_31_X23/X0/M3_g N_X23/7_X23/X0/M3_s
+ N_VDD_X23/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX23/X1/M0 N_X23/X1/6_X23/X1/M0_d N_STATE0_X23/X1/M0_g N_VSS_X23/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX23/X1/M1 N_X23/9_X23/X1/M1_d N_INIT2_X23/X1/M1_g N_X23/X1/6_X23/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX23/X1/M2 N_X23/9_X23/X1/M2_d N_STATE0_X23/X1/M2_g N_VDD_X23/X1/M2_s
+ N_VDD_X23/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX23/X1/M3 N_VDD_X23/X1/M3_d N_INIT2_X23/X1/M3_g N_X23/9_X23/X1/M3_s
+ N_VDD_X23/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX23/X2/M0 N_X23/X2/6_X23/X2/M0_d N_X23/9_X23/X2/M0_g N_VSS_X23/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX23/X2/M1 N_32_X23/X2/M1_d N_X23/7_X23/X2/M1_g N_X23/X2/6_X23/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX23/X2/M2 N_32_X23/X2/M2_d N_X23/9_X23/X2/M2_g N_VDD_X23/X2/M2_s
+ N_VDD_X23/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX23/X2/M3 N_VDD_X23/X2/M3_d N_X23/7_X23/X2/M3_g N_32_X23/X2/M3_s
+ N_VDD_X23/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX23/X3/M0 N_X23/8_X23/X3/M0_d N_STATE0_X23/X3/M0_g N_VSS_X23/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX23/X3/M1 N_X23/8_X23/X3/M1_d N_STATE0_X23/X3/M1_g N_VDD_X23/X3/M1_s
+ N_VDD_X23/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX24/X0/M0 N_X24/X0/6_X24/X0/M0_d N_X24/8_X24/X0/M0_g N_VSS_X24/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX24/X0/M1 N_X24/7_X24/X0/M1_d N_INIT2_X24/X0/M1_g N_X24/X0/6_X24/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX24/X0/M2 N_X24/7_X24/X0/M2_d N_X24/8_X24/X0/M2_g N_VDD_X24/X0/M2_s
+ N_VDD_X24/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX24/X0/M3 N_VDD_X24/X0/M3_d N_INIT2_X24/X0/M3_g N_X24/7_X24/X0/M3_s
+ N_VDD_X24/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX24/X1/M0 N_X24/X1/6_X24/X1/M0_d N_11_X24/X1/M0_g N_VSS_X24/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX24/X1/M1 N_X24/9_X24/X1/M1_d N_6_X24/X1/M1_g N_X24/X1/6_X24/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX24/X1/M2 N_X24/9_X24/X1/M2_d N_11_X24/X1/M2_g N_VDD_X24/X1/M2_s
+ N_VDD_X24/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX24/X1/M3 N_VDD_X24/X1/M3_d N_6_X24/X1/M3_g N_X24/9_X24/X1/M3_s
+ N_VDD_X24/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX24/X2/M0 N_X24/X2/6_X24/X2/M0_d N_X24/9_X24/X2/M0_g N_VSS_X24/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX24/X2/M1 N_33_X24/X2/M1_d N_X24/7_X24/X2/M1_g N_X24/X2/6_X24/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX24/X2/M2 N_33_X24/X2/M2_d N_X24/9_X24/X2/M2_g N_VDD_X24/X2/M2_s
+ N_VDD_X24/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX24/X2/M3 N_VDD_X24/X2/M3_d N_X24/7_X24/X2/M3_g N_33_X24/X2/M3_s
+ N_VDD_X24/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX24/X3/M0 N_X24/8_X24/X3/M0_d N_11_X24/X3/M0_g N_VSS_X24/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX24/X3/M1 N_X24/8_X24/X3/M1_d N_11_X24/X3/M1_g N_VDD_X24/X3/M1_s
+ N_VDD_X24/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX25/X0/M0 N_X25/X0/6_X25/X0/M0_d N_X25/8_X25/X0/M0_g N_VSS_X25/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX25/X0/M1 N_X25/7_X25/X0/M1_d N_35_X25/X0/M1_g N_X25/X0/6_X25/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX25/X0/M2 N_X25/7_X25/X0/M2_d N_X25/8_X25/X0/M2_g N_VDD_X25/X0/M2_s
+ N_VDD_X25/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX25/X0/M3 N_VDD_X25/X0/M3_d N_35_X25/X0/M3_g N_X25/7_X25/X0/M3_s
+ N_VDD_X25/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX25/X1/M0 N_X25/X1/6_X25/X1/M0_d N_STATE0_X25/X1/M0_g N_VSS_X25/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX25/X1/M1 N_X25/9_X25/X1/M1_d N_INIT3_X25/X1/M1_g N_X25/X1/6_X25/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX25/X1/M2 N_X25/9_X25/X1/M2_d N_STATE0_X25/X1/M2_g N_VDD_X25/X1/M2_s
+ N_VDD_X25/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX25/X1/M3 N_VDD_X25/X1/M3_d N_INIT3_X25/X1/M3_g N_X25/9_X25/X1/M3_s
+ N_VDD_X25/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX25/X2/M0 N_X25/X2/6_X25/X2/M0_d N_X25/9_X25/X2/M0_g N_VSS_X25/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX25/X2/M1 N_36_X25/X2/M1_d N_X25/7_X25/X2/M1_g N_X25/X2/6_X25/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX25/X2/M2 N_36_X25/X2/M2_d N_X25/9_X25/X2/M2_g N_VDD_X25/X2/M2_s
+ N_VDD_X25/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX25/X2/M3 N_VDD_X25/X2/M3_d N_X25/7_X25/X2/M3_g N_36_X25/X2/M3_s
+ N_VDD_X25/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX25/X3/M0 N_X25/8_X25/X3/M0_d N_STATE0_X25/X3/M0_g N_VSS_X25/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX25/X3/M1 N_X25/8_X25/X3/M1_d N_STATE0_X25/X3/M1_g N_VDD_X25/X3/M1_s
+ N_VDD_X25/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX26/X0/M0 N_X26/X0/6_X26/X0/M0_d N_X26/8_X26/X0/M0_g N_VSS_X26/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX26/X0/M1 N_X26/7_X26/X0/M1_d N_INIT3_X26/X0/M1_g N_X26/X0/6_X26/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX26/X0/M2 N_X26/7_X26/X0/M2_d N_X26/8_X26/X0/M2_g N_VDD_X26/X0/M2_s
+ N_VDD_X26/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX26/X0/M3 N_VDD_X26/X0/M3_d N_INIT3_X26/X0/M3_g N_X26/7_X26/X0/M3_s
+ N_VDD_X26/X0/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX26/X1/M0 N_X26/X1/6_X26/X1/M0_d N_11_X26/X1/M0_g N_VSS_X26/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX26/X1/M1 N_X26/9_X26/X1/M1_d N_8_X26/X1/M1_g N_X26/X1/6_X26/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX26/X1/M2 N_X26/9_X26/X1/M2_d N_11_X26/X1/M2_g N_VDD_X26/X1/M2_s
+ N_VDD_X26/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX26/X1/M3 N_VDD_X26/X1/M3_d N_8_X26/X1/M3_g N_X26/9_X26/X1/M3_s
+ N_VDD_X26/X1/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX26/X2/M0 N_X26/X2/6_X26/X2/M0_d N_X26/9_X26/X2/M0_g N_VSS_X26/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX26/X2/M1 N_37_X26/X2/M1_d N_X26/7_X26/X2/M1_g N_X26/X2/6_X26/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX26/X2/M2 N_37_X26/X2/M2_d N_X26/9_X26/X2/M2_g N_VDD_X26/X2/M2_s
+ N_VDD_X26/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX26/X2/M3 N_VDD_X26/X2/M3_d N_X26/7_X26/X2/M3_g N_37_X26/X2/M3_s
+ N_VDD_X26/X2/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX26/X3/M0 N_X26/8_X26/X3/M0_d N_11_X26/X3/M0_g N_VSS_X26/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=9.1e-13 PD=2.82e-06
+ PS=2.82e-06
mX26/X3/M1 N_X26/8_X26/X3/M1_d N_11_X26/X3/M1_g N_VDD_X26/X3/M1_s
+ N_VDD_X26/X3/M1_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=2.275e-12
+ PD=4.32e-06 PS=4.32e-06
mX27/X0/M0 N_X27/X0/11_X27/X0/M0_d N_X27/X0/7_X27/X0/M0_g N_VSS_X27/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX27/X0/M1 N_X27/X0/12_X27/X0/M1_d N_CLK_X27/X0/M1_g N_X27/X0/11_X27/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX27/X0/M2 N_X27/X0/9_X27/X0/M2_d N_X27/X0/8_X27/X0/M2_g N_X27/X0/12_X27/X0/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX27/X0/M3 N_X27/X0/9_X27/X0/M3_d N_X27/X0/7_X27/X0/M3_g N_VDD_X27/X0/M3_s
+ N_VDD_X27/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX27/X0/M4 N_VDD_X27/X0/M4_d N_CLK_X27/X0/M4_g N_X27/X0/9_X27/X0/M4_s
+ N_VDD_X27/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX27/X0/M5 N_X27/X0/9_X27/X0/M5_d N_X27/X0/8_X27/X0/M5_g N_VDD_X27/X0/M5_s
+ N_VDD_X27/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX27/X0/X6/M0 N_X27/X0/X6/6_X27/X0/X6/M0_d N_X27/X0/8_X27/X0/X6/M0_g
+ N_VSS_X27/X0/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X0/X6/M1 N_X27/X0/10_X27/X0/X6/M1_d N_X27/X0/7_X27/X0/X6/M1_g
+ N_X27/X0/X6/6_X27/X0/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X0/X6/M2 N_X27/X0/10_X27/X0/X6/M2_d N_X27/X0/8_X27/X0/X6/M2_g
+ N_VDD_X27/X0/X6/M2_s N_VDD_X27/X0/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X0/X6/M3 N_VDD_X27/X0/X6/M3_d N_X27/X0/7_X27/X0/X6/M3_g
+ N_X27/X0/10_X27/X0/X6/M3_s N_VDD_X27/X0/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X0/X7/M0 N_X27/X0/X7/6_X27/X0/X7/M0_d N_X27/X0/10_X27/X0/X7/M0_g
+ N_VSS_X27/X0/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X0/X7/M1 N_X27/X0/7_X27/X0/X7/M1_d N_CLK_X27/X0/X7/M1_g
+ N_X27/X0/X7/6_X27/X0/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X0/X7/M2 N_X27/X0/7_X27/X0/X7/M2_d N_X27/X0/10_X27/X0/X7/M2_g
+ N_VDD_X27/X0/X7/M2_s N_VDD_X27/X0/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X0/X7/M3 N_VDD_X27/X0/X7/M3_d N_CLK_X27/X0/X7/M3_g
+ N_X27/X0/7_X27/X0/X7/M3_s N_VDD_X27/X0/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X0/X8/M0 N_X27/X0/X8/6_X27/X0/X8/M0_d N_X27/X0/7_X27/X0/X8/M0_g
+ N_VSS_X27/X0/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X0/X8/M1 N_INIT0_X27/X0/X8/M1_d N_X27/12_X27/X0/X8/M1_g
+ N_X27/X0/X8/6_X27/X0/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X0/X8/M2 N_INIT0_X27/X0/X8/M2_d N_X27/X0/7_X27/X0/X8/M2_g
+ N_VDD_X27/X0/X8/M2_s N_VDD_X27/X0/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X0/X8/M3 N_VDD_X27/X0/X8/M3_d N_X27/12_X27/X0/X8/M3_g
+ N_INIT0_X27/X0/X8/M3_s N_VDD_X27/X0/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X0/X9/M0 N_X27/X0/X9/6_X27/X0/X9/M0_d N_INIT0_X27/X0/X9/M0_g
+ N_VSS_X27/X0/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X0/X9/M1 N_X27/12_X27/X0/X9/M1_d N_X27/X0/9_X27/X0/X9/M1_g
+ N_X27/X0/X9/6_X27/X0/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X0/X9/M2 N_X27/12_X27/X0/X9/M2_d N_INIT0_X27/X0/X9/M2_g
+ N_VDD_X27/X0/X9/M2_s N_VDD_X27/X0/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X0/X9/M3 N_VDD_X27/X0/X9/M3_d N_X27/X0/9_X27/X0/X9/M3_g
+ N_X27/12_X27/X0/X9/M3_s N_VDD_X27/X0/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X0/X10/M0 N_X27/X0/X10/6_X27/X0/X10/M0_d N_X27/X0/9_X27/X0/X10/M0_g
+ N_VSS_X27/X0/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X0/X10/M1 N_X27/X0/8_X27/X0/X10/M1_d N_17_X27/X0/X10/M1_g
+ N_X27/X0/X10/6_X27/X0/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X0/X10/M2 N_X27/X0/8_X27/X0/X10/M2_d N_X27/X0/9_X27/X0/X10/M2_g
+ N_VDD_X27/X0/X10/M2_s N_VDD_X27/X0/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X0/X10/M3 N_VDD_X27/X0/X10/M3_d N_17_X27/X0/X10/M3_g
+ N_X27/X0/8_X27/X0/X10/M3_s N_VDD_X27/X0/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X1/M0 N_X27/X1/11_X27/X1/M0_d N_X27/X1/7_X27/X1/M0_g N_VSS_X27/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX27/X1/M1 N_X27/X1/12_X27/X1/M1_d N_CLK_X27/X1/M1_g N_X27/X1/11_X27/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX27/X1/M2 N_X27/X1/9_X27/X1/M2_d N_X27/X1/8_X27/X1/M2_g N_X27/X1/12_X27/X1/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX27/X1/M3 N_X27/X1/9_X27/X1/M3_d N_X27/X1/7_X27/X1/M3_g N_VDD_X27/X1/M3_s
+ N_VDD_X27/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX27/X1/M4 N_VDD_X27/X1/M4_d N_CLK_X27/X1/M4_g N_X27/X1/9_X27/X1/M4_s
+ N_VDD_X27/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX27/X1/M5 N_X27/X1/9_X27/X1/M5_d N_X27/X1/8_X27/X1/M5_g N_VDD_X27/X1/M5_s
+ N_VDD_X27/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX27/X1/X6/M0 N_X27/X1/X6/6_X27/X1/X6/M0_d N_X27/X1/8_X27/X1/X6/M0_g
+ N_VSS_X27/X1/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X1/X6/M1 N_X27/X1/10_X27/X1/X6/M1_d N_X27/X1/7_X27/X1/X6/M1_g
+ N_X27/X1/X6/6_X27/X1/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X1/X6/M2 N_X27/X1/10_X27/X1/X6/M2_d N_X27/X1/8_X27/X1/X6/M2_g
+ N_VDD_X27/X1/X6/M2_s N_VDD_X27/X1/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X1/X6/M3 N_VDD_X27/X1/X6/M3_d N_X27/X1/7_X27/X1/X6/M3_g
+ N_X27/X1/10_X27/X1/X6/M3_s N_VDD_X27/X1/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X1/X7/M0 N_X27/X1/X7/6_X27/X1/X7/M0_d N_X27/X1/10_X27/X1/X7/M0_g
+ N_VSS_X27/X1/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X1/X7/M1 N_X27/X1/7_X27/X1/X7/M1_d N_CLK_X27/X1/X7/M1_g
+ N_X27/X1/X7/6_X27/X1/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X1/X7/M2 N_X27/X1/7_X27/X1/X7/M2_d N_X27/X1/10_X27/X1/X7/M2_g
+ N_VDD_X27/X1/X7/M2_s N_VDD_X27/X1/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X1/X7/M3 N_VDD_X27/X1/X7/M3_d N_CLK_X27/X1/X7/M3_g
+ N_X27/X1/7_X27/X1/X7/M3_s N_VDD_X27/X1/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X1/X8/M0 N_X27/X1/X8/6_X27/X1/X8/M0_d N_X27/X1/7_X27/X1/X8/M0_g
+ N_VSS_X27/X1/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X1/X8/M1 N_INIT1_X27/X1/X8/M1_d N_X27/13_X27/X1/X8/M1_g
+ N_X27/X1/X8/6_X27/X1/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X1/X8/M2 N_INIT1_X27/X1/X8/M2_d N_X27/X1/7_X27/X1/X8/M2_g
+ N_VDD_X27/X1/X8/M2_s N_VDD_X27/X1/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X1/X8/M3 N_VDD_X27/X1/X8/M3_d N_X27/13_X27/X1/X8/M3_g
+ N_INIT1_X27/X1/X8/M3_s N_VDD_X27/X1/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X1/X9/M0 N_X27/X1/X9/6_X27/X1/X9/M0_d N_INIT1_X27/X1/X9/M0_g
+ N_VSS_X27/X1/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X1/X9/M1 N_X27/13_X27/X1/X9/M1_d N_X27/X1/9_X27/X1/X9/M1_g
+ N_X27/X1/X9/6_X27/X1/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X1/X9/M2 N_X27/13_X27/X1/X9/M2_d N_INIT1_X27/X1/X9/M2_g
+ N_VDD_X27/X1/X9/M2_s N_VDD_X27/X1/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X1/X9/M3 N_VDD_X27/X1/X9/M3_d N_X27/X1/9_X27/X1/X9/M3_g
+ N_X27/13_X27/X1/X9/M3_s N_VDD_X27/X1/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X1/X10/M0 N_X27/X1/X10/6_X27/X1/X10/M0_d N_X27/X1/9_X27/X1/X10/M0_g
+ N_VSS_X27/X1/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X1/X10/M1 N_X27/X1/8_X27/X1/X10/M1_d N_27_X27/X1/X10/M1_g
+ N_X27/X1/X10/6_X27/X1/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X1/X10/M2 N_X27/X1/8_X27/X1/X10/M2_d N_X27/X1/9_X27/X1/X10/M2_g
+ N_VDD_X27/X1/X10/M2_s N_VDD_X27/X1/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X1/X10/M3 N_VDD_X27/X1/X10/M3_d N_27_X27/X1/X10/M3_g
+ N_X27/X1/8_X27/X1/X10/M3_s N_VDD_X27/X1/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X2/M0 N_X27/X2/11_X27/X2/M0_d N_X27/X2/7_X27/X2/M0_g N_VSS_X27/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX27/X2/M1 N_X27/X2/12_X27/X2/M1_d N_CLK_X27/X2/M1_g N_X27/X2/11_X27/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX27/X2/M2 N_X27/X2/9_X27/X2/M2_d N_X27/X2/8_X27/X2/M2_g N_X27/X2/12_X27/X2/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX27/X2/M3 N_X27/X2/9_X27/X2/M3_d N_X27/X2/7_X27/X2/M3_g N_VDD_X27/X2/M3_s
+ N_VDD_X27/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX27/X2/M4 N_VDD_X27/X2/M4_d N_CLK_X27/X2/M4_g N_X27/X2/9_X27/X2/M4_s
+ N_VDD_X27/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX27/X2/M5 N_X27/X2/9_X27/X2/M5_d N_X27/X2/8_X27/X2/M5_g N_VDD_X27/X2/M5_s
+ N_VDD_X27/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX27/X2/X6/M0 N_X27/X2/X6/6_X27/X2/X6/M0_d N_X27/X2/8_X27/X2/X6/M0_g
+ N_VSS_X27/X2/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X2/X6/M1 N_X27/X2/10_X27/X2/X6/M1_d N_X27/X2/7_X27/X2/X6/M1_g
+ N_X27/X2/X6/6_X27/X2/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X2/X6/M2 N_X27/X2/10_X27/X2/X6/M2_d N_X27/X2/8_X27/X2/X6/M2_g
+ N_VDD_X27/X2/X6/M2_s N_VDD_X27/X2/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X2/X6/M3 N_VDD_X27/X2/X6/M3_d N_X27/X2/7_X27/X2/X6/M3_g
+ N_X27/X2/10_X27/X2/X6/M3_s N_VDD_X27/X2/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X2/X7/M0 N_X27/X2/X7/6_X27/X2/X7/M0_d N_X27/X2/10_X27/X2/X7/M0_g
+ N_VSS_X27/X2/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X2/X7/M1 N_X27/X2/7_X27/X2/X7/M1_d N_CLK_X27/X2/X7/M1_g
+ N_X27/X2/X7/6_X27/X2/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X2/X7/M2 N_X27/X2/7_X27/X2/X7/M2_d N_X27/X2/10_X27/X2/X7/M2_g
+ N_VDD_X27/X2/X7/M2_s N_VDD_X27/X2/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X2/X7/M3 N_VDD_X27/X2/X7/M3_d N_CLK_X27/X2/X7/M3_g
+ N_X27/X2/7_X27/X2/X7/M3_s N_VDD_X27/X2/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X2/X8/M0 N_X27/X2/X8/6_X27/X2/X8/M0_d N_X27/X2/7_X27/X2/X8/M0_g
+ N_VSS_X27/X2/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X2/X8/M1 N_INIT2_X27/X2/X8/M1_d N_X27/14_X27/X2/X8/M1_g
+ N_X27/X2/X8/6_X27/X2/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X2/X8/M2 N_INIT2_X27/X2/X8/M2_d N_X27/X2/7_X27/X2/X8/M2_g
+ N_VDD_X27/X2/X8/M2_s N_VDD_X27/X2/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X2/X8/M3 N_VDD_X27/X2/X8/M3_d N_X27/14_X27/X2/X8/M3_g
+ N_INIT2_X27/X2/X8/M3_s N_VDD_X27/X2/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X2/X9/M0 N_X27/X2/X9/6_X27/X2/X9/M0_d N_INIT2_X27/X2/X9/M0_g
+ N_VSS_X27/X2/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X2/X9/M1 N_X27/14_X27/X2/X9/M1_d N_X27/X2/9_X27/X2/X9/M1_g
+ N_X27/X2/X9/6_X27/X2/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X2/X9/M2 N_X27/14_X27/X2/X9/M2_d N_INIT2_X27/X2/X9/M2_g
+ N_VDD_X27/X2/X9/M2_s N_VDD_X27/X2/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X2/X9/M3 N_VDD_X27/X2/X9/M3_d N_X27/X2/9_X27/X2/X9/M3_g
+ N_X27/14_X27/X2/X9/M3_s N_VDD_X27/X2/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X2/X10/M0 N_X27/X2/X10/6_X27/X2/X10/M0_d N_X27/X2/9_X27/X2/X10/M0_g
+ N_VSS_X27/X2/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X2/X10/M1 N_X27/X2/8_X27/X2/X10/M1_d N_33_X27/X2/X10/M1_g
+ N_X27/X2/X10/6_X27/X2/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X2/X10/M2 N_X27/X2/8_X27/X2/X10/M2_d N_X27/X2/9_X27/X2/X10/M2_g
+ N_VDD_X27/X2/X10/M2_s N_VDD_X27/X2/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X2/X10/M3 N_VDD_X27/X2/X10/M3_d N_33_X27/X2/X10/M3_g
+ N_X27/X2/8_X27/X2/X10/M3_s N_VDD_X27/X2/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X3/M0 N_X27/X3/11_X27/X3/M0_d N_X27/X3/7_X27/X3/M0_g N_VSS_X27/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX27/X3/M1 N_X27/X3/12_X27/X3/M1_d N_CLK_X27/X3/M1_g N_X27/X3/11_X27/X3/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX27/X3/M2 N_X27/X3/9_X27/X3/M2_d N_X27/X3/8_X27/X3/M2_g N_X27/X3/12_X27/X3/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX27/X3/M3 N_X27/X3/9_X27/X3/M3_d N_X27/X3/7_X27/X3/M3_g N_VDD_X27/X3/M3_s
+ N_VDD_X27/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX27/X3/M4 N_VDD_X27/X3/M4_d N_CLK_X27/X3/M4_g N_X27/X3/9_X27/X3/M4_s
+ N_VDD_X27/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX27/X3/M5 N_X27/X3/9_X27/X3/M5_d N_X27/X3/8_X27/X3/M5_g N_VDD_X27/X3/M5_s
+ N_VDD_X27/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX27/X3/X6/M0 N_X27/X3/X6/6_X27/X3/X6/M0_d N_X27/X3/8_X27/X3/X6/M0_g
+ N_VSS_X27/X3/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X3/X6/M1 N_X27/X3/10_X27/X3/X6/M1_d N_X27/X3/7_X27/X3/X6/M1_g
+ N_X27/X3/X6/6_X27/X3/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X3/X6/M2 N_X27/X3/10_X27/X3/X6/M2_d N_X27/X3/8_X27/X3/X6/M2_g
+ N_VDD_X27/X3/X6/M2_s N_VDD_X27/X3/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X3/X6/M3 N_VDD_X27/X3/X6/M3_d N_X27/X3/7_X27/X3/X6/M3_g
+ N_X27/X3/10_X27/X3/X6/M3_s N_VDD_X27/X3/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X3/X7/M0 N_X27/X3/X7/6_X27/X3/X7/M0_d N_X27/X3/10_X27/X3/X7/M0_g
+ N_VSS_X27/X3/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X3/X7/M1 N_X27/X3/7_X27/X3/X7/M1_d N_CLK_X27/X3/X7/M1_g
+ N_X27/X3/X7/6_X27/X3/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X3/X7/M2 N_X27/X3/7_X27/X3/X7/M2_d N_X27/X3/10_X27/X3/X7/M2_g
+ N_VDD_X27/X3/X7/M2_s N_VDD_X27/X3/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X3/X7/M3 N_VDD_X27/X3/X7/M3_d N_CLK_X27/X3/X7/M3_g
+ N_X27/X3/7_X27/X3/X7/M3_s N_VDD_X27/X3/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X3/X8/M0 N_X27/X3/X8/6_X27/X3/X8/M0_d N_X27/X3/7_X27/X3/X8/M0_g
+ N_VSS_X27/X3/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X3/X8/M1 N_INIT3_X27/X3/X8/M1_d N_X27/15_X27/X3/X8/M1_g
+ N_X27/X3/X8/6_X27/X3/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X3/X8/M2 N_INIT3_X27/X3/X8/M2_d N_X27/X3/7_X27/X3/X8/M2_g
+ N_VDD_X27/X3/X8/M2_s N_VDD_X27/X3/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X3/X8/M3 N_VDD_X27/X3/X8/M3_d N_X27/15_X27/X3/X8/M3_g
+ N_INIT3_X27/X3/X8/M3_s N_VDD_X27/X3/X8/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X3/X9/M0 N_X27/X3/X9/6_X27/X3/X9/M0_d N_INIT3_X27/X3/X9/M0_g
+ N_VSS_X27/X3/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X3/X9/M1 N_X27/15_X27/X3/X9/M1_d N_X27/X3/9_X27/X3/X9/M1_g
+ N_X27/X3/X9/6_X27/X3/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X3/X9/M2 N_X27/15_X27/X3/X9/M2_d N_INIT3_X27/X3/X9/M2_g
+ N_VDD_X27/X3/X9/M2_s N_VDD_X27/X3/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X3/X9/M3 N_VDD_X27/X3/X9/M3_d N_X27/X3/9_X27/X3/X9/M3_g
+ N_X27/15_X27/X3/X9/M3_s N_VDD_X27/X3/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX27/X3/X10/M0 N_X27/X3/X10/6_X27/X3/X10/M0_d N_X27/X3/9_X27/X3/X10/M0_g
+ N_VSS_X27/X3/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX27/X3/X10/M1 N_X27/X3/8_X27/X3/X10/M1_d N_37_X27/X3/X10/M1_g
+ N_X27/X3/X10/6_X27/X3/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX27/X3/X10/M2 N_X27/X3/8_X27/X3/X10/M2_d N_X27/X3/9_X27/X3/X10/M2_g
+ N_VDD_X27/X3/X10/M2_s N_VDD_X27/X3/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX27/X3/X10/M3 N_VDD_X27/X3/X10/M3_d N_37_X27/X3/X10/M3_g
+ N_X27/X3/8_X27/X3/X10/M3_s N_VDD_X27/X3/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X0/M0 N_X28/X0/11_X28/X0/M0_d N_X28/X0/7_X28/X0/M0_g N_VSS_X28/X0/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX28/X0/M1 N_X28/X0/12_X28/X0/M1_d N_CLK_X28/X0/M1_g N_X28/X0/11_X28/X0/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX28/X0/M2 N_X28/X0/9_X28/X0/M2_d N_X28/X0/8_X28/X0/M2_g N_X28/X0/12_X28/X0/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX28/X0/M3 N_X28/X0/9_X28/X0/M3_d N_X28/X0/7_X28/X0/M3_g N_VDD_X28/X0/M3_s
+ N_VDD_X28/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X0/M4 N_VDD_X28/X0/M4_d N_CLK_X28/X0/M4_g N_X28/X0/9_X28/X0/M4_s
+ N_VDD_X28/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX28/X0/M5 N_X28/X0/9_X28/X0/M5_d N_X28/X0/8_X28/X0/M5_g N_VDD_X28/X0/M5_s
+ N_VDD_X28/X0/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X0/X6/M0 N_X28/X0/X6/6_X28/X0/X6/M0_d N_X28/X0/8_X28/X0/X6/M0_g
+ N_VSS_X28/X0/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X0/X6/M1 N_X28/X0/10_X28/X0/X6/M1_d N_X28/X0/7_X28/X0/X6/M1_g
+ N_X28/X0/X6/6_X28/X0/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X0/X6/M2 N_X28/X0/10_X28/X0/X6/M2_d N_X28/X0/8_X28/X0/X6/M2_g
+ N_VDD_X28/X0/X6/M2_s N_VDD_X28/X0/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X0/X6/M3 N_VDD_X28/X0/X6/M3_d N_X28/X0/7_X28/X0/X6/M3_g
+ N_X28/X0/10_X28/X0/X6/M3_s N_VDD_X28/X0/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X0/X7/M0 N_X28/X0/X7/6_X28/X0/X7/M0_d N_X28/X0/10_X28/X0/X7/M0_g
+ N_VSS_X28/X0/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X0/X7/M1 N_X28/X0/7_X28/X0/X7/M1_d N_CLK_X28/X0/X7/M1_g
+ N_X28/X0/X7/6_X28/X0/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X0/X7/M2 N_X28/X0/7_X28/X0/X7/M2_d N_X28/X0/10_X28/X0/X7/M2_g
+ N_VDD_X28/X0/X7/M2_s N_VDD_X28/X0/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X0/X7/M3 N_VDD_X28/X0/X7/M3_d N_CLK_X28/X0/X7/M3_g
+ N_X28/X0/7_X28/X0/X7/M3_s N_VDD_X28/X0/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X0/X8/M0 N_X28/X0/X8/6_X28/X0/X8/M0_d N_X28/X0/7_X28/X0/X8/M0_g
+ N_VSS_X28/X0/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X0/X8/M1 N_12_X28/X0/X8/M1_d N_X28/12_X28/X0/X8/M1_g
+ N_X28/X0/X8/6_X28/X0/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X0/X8/M2 N_12_X28/X0/X8/M2_d N_X28/X0/7_X28/X0/X8/M2_g N_VDD_X28/X0/X8/M2_s
+ N_VDD_X28/X0/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X0/X8/M3 N_VDD_X28/X0/X8/M3_d N_X28/12_X28/X0/X8/M3_g N_12_X28/X0/X8/M3_s
+ N_VDD_X28/X0/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X0/X9/M0 N_X28/X0/X9/6_X28/X0/X9/M0_d N_12_X28/X0/X9/M0_g
+ N_VSS_X28/X0/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X0/X9/M1 N_X28/12_X28/X0/X9/M1_d N_X28/X0/9_X28/X0/X9/M1_g
+ N_X28/X0/X9/6_X28/X0/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X0/X9/M2 N_X28/12_X28/X0/X9/M2_d N_12_X28/X0/X9/M2_g N_VDD_X28/X0/X9/M2_s
+ N_VDD_X28/X0/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X0/X9/M3 N_VDD_X28/X0/X9/M3_d N_X28/X0/9_X28/X0/X9/M3_g
+ N_X28/12_X28/X0/X9/M3_s N_VDD_X28/X0/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X0/X10/M0 N_X28/X0/X10/6_X28/X0/X10/M0_d N_X28/X0/9_X28/X0/X10/M0_g
+ N_VSS_X28/X0/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X0/X10/M1 N_X28/X0/8_X28/X0/X10/M1_d N_M0_X28/X0/X10/M1_g
+ N_X28/X0/X10/6_X28/X0/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X0/X10/M2 N_X28/X0/8_X28/X0/X10/M2_d N_X28/X0/9_X28/X0/X10/M2_g
+ N_VDD_X28/X0/X10/M2_s N_VDD_X28/X0/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X0/X10/M3 N_VDD_X28/X0/X10/M3_d N_M0_X28/X0/X10/M3_g
+ N_X28/X0/8_X28/X0/X10/M3_s N_VDD_X28/X0/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X1/M0 N_X28/X1/11_X28/X1/M0_d N_X28/X1/7_X28/X1/M0_g N_VSS_X28/X1/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX28/X1/M1 N_X28/X1/12_X28/X1/M1_d N_CLK_X28/X1/M1_g N_X28/X1/11_X28/X1/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX28/X1/M2 N_X28/X1/9_X28/X1/M2_d N_X28/X1/8_X28/X1/M2_g N_X28/X1/12_X28/X1/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX28/X1/M3 N_X28/X1/9_X28/X1/M3_d N_X28/X1/7_X28/X1/M3_g N_VDD_X28/X1/M3_s
+ N_VDD_X28/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X1/M4 N_VDD_X28/X1/M4_d N_CLK_X28/X1/M4_g N_X28/X1/9_X28/X1/M4_s
+ N_VDD_X28/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX28/X1/M5 N_X28/X1/9_X28/X1/M5_d N_X28/X1/8_X28/X1/M5_g N_VDD_X28/X1/M5_s
+ N_VDD_X28/X1/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X1/X6/M0 N_X28/X1/X6/6_X28/X1/X6/M0_d N_X28/X1/8_X28/X1/X6/M0_g
+ N_VSS_X28/X1/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X1/X6/M1 N_X28/X1/10_X28/X1/X6/M1_d N_X28/X1/7_X28/X1/X6/M1_g
+ N_X28/X1/X6/6_X28/X1/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X1/X6/M2 N_X28/X1/10_X28/X1/X6/M2_d N_X28/X1/8_X28/X1/X6/M2_g
+ N_VDD_X28/X1/X6/M2_s N_VDD_X28/X1/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X1/X6/M3 N_VDD_X28/X1/X6/M3_d N_X28/X1/7_X28/X1/X6/M3_g
+ N_X28/X1/10_X28/X1/X6/M3_s N_VDD_X28/X1/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X1/X7/M0 N_X28/X1/X7/6_X28/X1/X7/M0_d N_X28/X1/10_X28/X1/X7/M0_g
+ N_VSS_X28/X1/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X1/X7/M1 N_X28/X1/7_X28/X1/X7/M1_d N_CLK_X28/X1/X7/M1_g
+ N_X28/X1/X7/6_X28/X1/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X1/X7/M2 N_X28/X1/7_X28/X1/X7/M2_d N_X28/X1/10_X28/X1/X7/M2_g
+ N_VDD_X28/X1/X7/M2_s N_VDD_X28/X1/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X1/X7/M3 N_VDD_X28/X1/X7/M3_d N_CLK_X28/X1/X7/M3_g
+ N_X28/X1/7_X28/X1/X7/M3_s N_VDD_X28/X1/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X1/X8/M0 N_X28/X1/X8/6_X28/X1/X8/M0_d N_X28/X1/7_X28/X1/X8/M0_g
+ N_VSS_X28/X1/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X1/X8/M1 N_24_X28/X1/X8/M1_d N_X28/13_X28/X1/X8/M1_g
+ N_X28/X1/X8/6_X28/X1/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X1/X8/M2 N_24_X28/X1/X8/M2_d N_X28/X1/7_X28/X1/X8/M2_g N_VDD_X28/X1/X8/M2_s
+ N_VDD_X28/X1/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X1/X8/M3 N_VDD_X28/X1/X8/M3_d N_X28/13_X28/X1/X8/M3_g N_24_X28/X1/X8/M3_s
+ N_VDD_X28/X1/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X1/X9/M0 N_X28/X1/X9/6_X28/X1/X9/M0_d N_24_X28/X1/X9/M0_g
+ N_VSS_X28/X1/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X1/X9/M1 N_X28/13_X28/X1/X9/M1_d N_X28/X1/9_X28/X1/X9/M1_g
+ N_X28/X1/X9/6_X28/X1/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X1/X9/M2 N_X28/13_X28/X1/X9/M2_d N_24_X28/X1/X9/M2_g N_VDD_X28/X1/X9/M2_s
+ N_VDD_X28/X1/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X1/X9/M3 N_VDD_X28/X1/X9/M3_d N_X28/X1/9_X28/X1/X9/M3_g
+ N_X28/13_X28/X1/X9/M3_s N_VDD_X28/X1/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X1/X10/M0 N_X28/X1/X10/6_X28/X1/X10/M0_d N_X28/X1/9_X28/X1/X10/M0_g
+ N_VSS_X28/X1/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X1/X10/M1 N_X28/X1/8_X28/X1/X10/M1_d N_M1_X28/X1/X10/M1_g
+ N_X28/X1/X10/6_X28/X1/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X1/X10/M2 N_X28/X1/8_X28/X1/X10/M2_d N_X28/X1/9_X28/X1/X10/M2_g
+ N_VDD_X28/X1/X10/M2_s N_VDD_X28/X1/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X1/X10/M3 N_VDD_X28/X1/X10/M3_d N_M1_X28/X1/X10/M3_g
+ N_X28/X1/8_X28/X1/X10/M3_s N_VDD_X28/X1/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X2/M0 N_X28/X2/11_X28/X2/M0_d N_X28/X2/7_X28/X2/M0_g N_VSS_X28/X2/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX28/X2/M1 N_X28/X2/12_X28/X2/M1_d N_CLK_X28/X2/M1_g N_X28/X2/11_X28/X2/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX28/X2/M2 N_X28/X2/9_X28/X2/M2_d N_X28/X2/8_X28/X2/M2_g N_X28/X2/12_X28/X2/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX28/X2/M3 N_X28/X2/9_X28/X2/M3_d N_X28/X2/7_X28/X2/M3_g N_VDD_X28/X2/M3_s
+ N_VDD_X28/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X2/M4 N_VDD_X28/X2/M4_d N_CLK_X28/X2/M4_g N_X28/X2/9_X28/X2/M4_s
+ N_VDD_X28/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX28/X2/M5 N_X28/X2/9_X28/X2/M5_d N_X28/X2/8_X28/X2/M5_g N_VDD_X28/X2/M5_s
+ N_VDD_X28/X2/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X2/X6/M0 N_X28/X2/X6/6_X28/X2/X6/M0_d N_X28/X2/8_X28/X2/X6/M0_g
+ N_VSS_X28/X2/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X2/X6/M1 N_X28/X2/10_X28/X2/X6/M1_d N_X28/X2/7_X28/X2/X6/M1_g
+ N_X28/X2/X6/6_X28/X2/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X2/X6/M2 N_X28/X2/10_X28/X2/X6/M2_d N_X28/X2/8_X28/X2/X6/M2_g
+ N_VDD_X28/X2/X6/M2_s N_VDD_X28/X2/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X2/X6/M3 N_VDD_X28/X2/X6/M3_d N_X28/X2/7_X28/X2/X6/M3_g
+ N_X28/X2/10_X28/X2/X6/M3_s N_VDD_X28/X2/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X2/X7/M0 N_X28/X2/X7/6_X28/X2/X7/M0_d N_X28/X2/10_X28/X2/X7/M0_g
+ N_VSS_X28/X2/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X2/X7/M1 N_X28/X2/7_X28/X2/X7/M1_d N_CLK_X28/X2/X7/M1_g
+ N_X28/X2/X7/6_X28/X2/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X2/X7/M2 N_X28/X2/7_X28/X2/X7/M2_d N_X28/X2/10_X28/X2/X7/M2_g
+ N_VDD_X28/X2/X7/M2_s N_VDD_X28/X2/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X2/X7/M3 N_VDD_X28/X2/X7/M3_d N_CLK_X28/X2/X7/M3_g
+ N_X28/X2/7_X28/X2/X7/M3_s N_VDD_X28/X2/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X2/X8/M0 N_X28/X2/X8/6_X28/X2/X8/M0_d N_X28/X2/7_X28/X2/X8/M0_g
+ N_VSS_X28/X2/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X2/X8/M1 N_31_X28/X2/X8/M1_d N_X28/14_X28/X2/X8/M1_g
+ N_X28/X2/X8/6_X28/X2/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X2/X8/M2 N_31_X28/X2/X8/M2_d N_X28/X2/7_X28/X2/X8/M2_g N_VDD_X28/X2/X8/M2_s
+ N_VDD_X28/X2/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X2/X8/M3 N_VDD_X28/X2/X8/M3_d N_X28/14_X28/X2/X8/M3_g N_31_X28/X2/X8/M3_s
+ N_VDD_X28/X2/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X2/X9/M0 N_X28/X2/X9/6_X28/X2/X9/M0_d N_31_X28/X2/X9/M0_g
+ N_VSS_X28/X2/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X2/X9/M1 N_X28/14_X28/X2/X9/M1_d N_X28/X2/9_X28/X2/X9/M1_g
+ N_X28/X2/X9/6_X28/X2/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X2/X9/M2 N_X28/14_X28/X2/X9/M2_d N_31_X28/X2/X9/M2_g N_VDD_X28/X2/X9/M2_s
+ N_VDD_X28/X2/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X2/X9/M3 N_VDD_X28/X2/X9/M3_d N_X28/X2/9_X28/X2/X9/M3_g
+ N_X28/14_X28/X2/X9/M3_s N_VDD_X28/X2/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X2/X10/M0 N_X28/X2/X10/6_X28/X2/X10/M0_d N_X28/X2/9_X28/X2/X10/M0_g
+ N_VSS_X28/X2/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X2/X10/M1 N_X28/X2/8_X28/X2/X10/M1_d N_M2_X28/X2/X10/M1_g
+ N_X28/X2/X10/6_X28/X2/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X2/X10/M2 N_X28/X2/8_X28/X2/X10/M2_d N_X28/X2/9_X28/X2/X10/M2_g
+ N_VDD_X28/X2/X10/M2_s N_VDD_X28/X2/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X2/X10/M3 N_VDD_X28/X2/X10/M3_d N_M2_X28/X2/X10/M3_g
+ N_X28/X2/8_X28/X2/X10/M3_s N_VDD_X28/X2/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X3/M0 N_X28/X3/11_X28/X3/M0_d N_X28/X3/7_X28/X3/M0_g N_VSS_X28/X3/M0_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=9.1e-13 PD=8.2e-07
+ PS=2.82e-06
mX28/X3/M1 N_X28/X3/12_X28/X3/M1_d N_CLK_X28/X3/M1_g N_X28/X3/11_X28/X3/M1_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13 AS=4.1e-13 PD=8.2e-07
+ PS=8.2e-07
mX28/X3/M2 N_X28/X3/9_X28/X3/M2_d N_X28/X3/8_X28/X3/M2_g N_X28/X3/12_X28/X3/M2_s
+ N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=9.1e-13 AS=4.1e-13 PD=2.82e-06
+ PS=8.2e-07
mX28/X3/M3 N_X28/X3/9_X28/X3/M3_d N_X28/X3/7_X28/X3/M3_g N_VDD_X28/X3/M3_s
+ N_VDD_X28/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X3/M4 N_VDD_X28/X3/M4_d N_CLK_X28/X3/M4_g N_X28/X3/9_X28/X3/M4_s
+ N_VDD_X28/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=1.025e-12
+ PD=8.2e-07 PS=8.2e-07
mX28/X3/M5 N_X28/X3/9_X28/X3/M5_d N_X28/X3/8_X28/X3/M5_g N_VDD_X28/X3/M5_s
+ N_VDD_X28/X3/M3_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X3/X6/M0 N_X28/X3/X6/6_X28/X3/X6/M0_d N_X28/X3/8_X28/X3/X6/M0_g
+ N_VSS_X28/X3/X6/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X3/X6/M1 N_X28/X3/10_X28/X3/X6/M1_d N_X28/X3/7_X28/X3/X6/M1_g
+ N_X28/X3/X6/6_X28/X3/X6/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X3/X6/M2 N_X28/X3/10_X28/X3/X6/M2_d N_X28/X3/8_X28/X3/X6/M2_g
+ N_VDD_X28/X3/X6/M2_s N_VDD_X28/X3/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X3/X6/M3 N_VDD_X28/X3/X6/M3_d N_X28/X3/7_X28/X3/X6/M3_g
+ N_X28/X3/10_X28/X3/X6/M3_s N_VDD_X28/X3/X6/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X3/X7/M0 N_X28/X3/X7/6_X28/X3/X7/M0_d N_X28/X3/10_X28/X3/X7/M0_g
+ N_VSS_X28/X3/X7/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X3/X7/M1 N_X28/X3/7_X28/X3/X7/M1_d N_CLK_X28/X3/X7/M1_g
+ N_X28/X3/X7/6_X28/X3/X7/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X3/X7/M2 N_X28/X3/7_X28/X3/X7/M2_d N_X28/X3/10_X28/X3/X7/M2_g
+ N_VDD_X28/X3/X7/M2_s N_VDD_X28/X3/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X3/X7/M3 N_VDD_X28/X3/X7/M3_d N_CLK_X28/X3/X7/M3_g
+ N_X28/X3/7_X28/X3/X7/M3_s N_VDD_X28/X3/X7/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X3/X8/M0 N_X28/X3/X8/6_X28/X3/X8/M0_d N_X28/X3/7_X28/X3/X8/M0_g
+ N_VSS_X28/X3/X8/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X3/X8/M1 N_35_X28/X3/X8/M1_d N_X28/15_X28/X3/X8/M1_g
+ N_X28/X3/X8/6_X28/X3/X8/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X3/X8/M2 N_35_X28/X3/X8/M2_d N_X28/X3/7_X28/X3/X8/M2_g N_VDD_X28/X3/X8/M2_s
+ N_VDD_X28/X3/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X3/X8/M3 N_VDD_X28/X3/X8/M3_d N_X28/15_X28/X3/X8/M3_g N_35_X28/X3/X8/M3_s
+ N_VDD_X28/X3/X8/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=2.275e-12 AS=1.025e-12
+ PD=4.32e-06 PS=8.2e-07
mX28/X3/X9/M0 N_X28/X3/X9/6_X28/X3/X9/M0_d N_35_X28/X3/X9/M0_g
+ N_VSS_X28/X3/X9/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X3/X9/M1 N_X28/15_X28/X3/X9/M1_d N_X28/X3/9_X28/X3/X9/M1_g
+ N_X28/X3/X9/6_X28/X3/X9/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X3/X9/M2 N_X28/15_X28/X3/X9/M2_d N_35_X28/X3/X9/M2_g N_VDD_X28/X3/X9/M2_s
+ N_VDD_X28/X3/X9/M2_b P_18 L=1.8e-07 W=2.5e-06 AD=1.025e-12 AS=2.275e-12
+ PD=8.2e-07 PS=4.32e-06
mX28/X3/X9/M3 N_VDD_X28/X3/X9/M3_d N_X28/X3/9_X28/X3/X9/M3_g
+ N_X28/15_X28/X3/X9/M3_s N_VDD_X28/X3/X9/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
mX28/X3/X10/M0 N_X28/X3/X10/6_X28/X3/X10/M0_d N_X28/X3/9_X28/X3/X10/M0_g
+ N_VSS_X28/X3/X10/M0_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06 AD=4.1e-13
+ AS=9.1e-13 PD=8.2e-07 PS=2.82e-06
mX28/X3/X10/M1 N_X28/X3/8_X28/X3/X10/M1_d N_M3_X28/X3/X10/M1_g
+ N_X28/X3/X10/6_X28/X3/X10/M1_s N_VSS_X0/X0/M0_b N_18 L=1.8e-07 W=1e-06
+ AD=9.1e-13 AS=4.1e-13 PD=2.82e-06 PS=8.2e-07
mX28/X3/X10/M2 N_X28/X3/8_X28/X3/X10/M2_d N_X28/X3/9_X28/X3/X10/M2_g
+ N_VDD_X28/X3/X10/M2_s N_VDD_X28/X3/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=1.025e-12 AS=2.275e-12 PD=8.2e-07 PS=4.32e-06
mX28/X3/X10/M3 N_VDD_X28/X3/X10/M3_d N_M3_X28/X3/X10/M3_g
+ N_X28/X3/8_X28/X3/X10/M3_s N_VDD_X28/X3/X10/M2_b P_18 L=1.8e-07 W=2.5e-06
+ AD=2.275e-12 AS=1.025e-12 PD=4.32e-06 PS=8.2e-07
*
.include "Coin_bank.pex.sp.COIN_BANK.pxi"
*
.ends
*
*
